`include "i2c_uvc/i2c_common.svh"
`include "i2c_uvc/i2c_transaction.svh"
`include "i2c_uvc/i2c_config.svh"
`include "i2c_uvc/i2c_adapter.svh"
`include "i2c_uvc/i2c_sequencer.svh"
`include "i2c_uvc/i2c_driver.svh"
`include "i2c_uvc/i2c_monitor.svh"
`include "i2c_uvc/i2c_agent.svh"
`include "i2c_uvc/i2c_sequence.svh"
