typedef class rcc_config;
typedef class rcc_driver;

`include "rcc_uvc/rcc_config.svh"
`include "rcc_uvc/rcc_driver.svh"
