
//------------------------------------------------------------------------------
// PACKAGE: tb_pkg
//
// Package for test bench
//------------------------------------------------------------------------------
package tb_pkg;
  `include "uvm_macros.svh"
  import uvm_pkg::*;
  import uvc_pkg::*;
  
  `include "tb_env.svh"
endpackage
