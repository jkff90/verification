typedef class amba_axi4_transaction;
typedef class amba_axi4_config;
typedef class amba_axi4_adapter;
typedef class amba_axi4_sequencer;
typedef class amba_axi4_driver;
typedef class amba_axi4_monitor;
typedef class amba_axi4_coverage;
typedef class amba_axi4_agent;
typedef class amba_axi4_pipelined_sequence;
typedef class amba_axi4_unpipelined_sequence;
typedef class amba_axi4_passthru_sequence;

`include "amba_axi4_uvc/amba_axi4_common.svh"
`include "amba_axi4_uvc/amba_axi4_transaction.svh"
`include "amba_axi4_uvc/amba_axi4_config.svh"
`include "amba_axi4_uvc/amba_axi4_adapter.svh"
`include "amba_axi4_uvc/amba_axi4_sequencer.svh"
`include "amba_axi4_uvc/amba_axi4_driver.svh"
`include "amba_axi4_uvc/amba_axi4_monitor.svh"
`include "amba_axi4_uvc/amba_axi4_coverage.svh"
`include "amba_axi4_uvc/amba_axi4_passive_device.svh"
`include "amba_axi4_uvc/amba_axi4_agent.svh"
`include "amba_axi4_uvc/amba_axi4_pipelined_sequence.svh"
`include "amba_axi4_uvc/amba_axi4_unpipelined_sequence.svh"
`include "amba_axi4_uvc/amba_axi4_passthru_sequence.svh"
