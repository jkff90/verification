`include "irq_uvc/irq_common.svh"
`include "irq_uvc/irq_transaction.svh"
`include "irq_uvc/irq_config.svh"
`include "irq_uvc/irq_adapter.svh"
`include "irq_uvc/irq_sequencer.svh"
`include "irq_uvc/irq_driver.svh"
`include "irq_uvc/irq_monitor.svh"
`include "irq_uvc/irq_agent.svh"
`include "irq_uvc/irq_sequence.svh"
