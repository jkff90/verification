
//------------------------------------------------------------------------------
// PACKAGE: toolbox
//
// Contains many useful tools for SystemVerilog programming
//------------------------------------------------------------------------------
package toolbox_pkg;
  `include "packages/toolbox/a2e.svh"
  `include "packages/toolbox/process_db.svh"
endpackage
