
`include "video_uvc/video_common.svh"
`include "video_uvc/video_transaction.svh"
`include "video_uvc/video_config.svh"
`include "video_uvc/video_adapter.svh"
`include "video_uvc/video_sequencer.svh"
`include "video_uvc/video_driver.svh"
`include "video_uvc/video_monitor.svh"
`include "video_uvc/video_recorder.svh"
`include "video_uvc/video_agent.svh"
`include "video_uvc/video_sequence.svh"
