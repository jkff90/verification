`include "avlmm_uvc/avlmm_common.svh"
`include "avlmm_uvc/avlmm_transaction.svh"
`include "avlmm_uvc/avlmm_config.svh"
`include "avlmm_uvc/avlmm_adapter.svh"
`include "avlmm_uvc/avlmm_sequencer.svh"
`include "avlmm_uvc/avlmm_driver.svh"
`include "avlmm_uvc/avlmm_monitor.svh"
`include "avlmm_uvc/avlmm_agent.svh"
`include "avlmm_uvc/avlmm_sequence.svh"
