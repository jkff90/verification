`include "reg_adapter_uvc/reg_adapter_wishbone.svh"
