
`include "scb_uvc/scb_config.svh"
`include "scb_uvc/two_sides_scb.svh"
