`include "adapter_uvc/adapter_base.svh"
`include "adapter_uvc/packet_to_avlst_adapter.svh"
`include "adapter_uvc/video_to_packet_adapter.svh"
