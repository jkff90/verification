
//------------------------------------------------------------------------------
// Package: sequence_pkg
//------------------------------------------------------------------------------
package sequence_pkg;
  `include "uvm_macros.svh"
  import uvm_pkg::*;
  import uvc_pkg::*;
  import tb_pkg::*;
  
  `include "sequence/dut_config_sequence.svh"
  `include "sequence/video_file_sequence.svh"
endpackage : sequence_pkg
