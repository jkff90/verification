//------------------------------------------------------------------------------
// Author: anonymous
// Email: anonymous@noreply.com
//------------------------------------------------------------------------------

//------------------------------------------------------------------------------
// Package: uvc_pkg
//
// UVM Verification Components package
//------------------------------------------------------------------------------
package uvc_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"
  
  `include "uvc.svh"
endpackage : uvc_pkg
