`include "amba_axi4_uvc/amba_axi4_uvc.svh"
`include "avlmm_uvc/avlmm_uvc.svh"
`include "avlst_uvc/avlst_uvc.svh"
`include "avlst_uvc/avlst_uvc.svh"
`include "i2c_uvc/i2c_uvc.svh"
`include "irq_uvc/irq_uvc.svh"
`include "packet_uvc/packet_uvc.svh"
`include "video_uvc/video_uvc.svh"
`include "wishbone_uvc/wishbone_uvc.svh"
`include "reg_adapter_uvc/reg_adapter_uvc.svh"
`include "adapter_uvc/adapter_uvc.svh"
`include "scb_uvc/scb_uvc.svh"
`include "env_uvc/env_uvc.svh"
