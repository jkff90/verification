`include "interfaces/backdoor_if.sv"
`include "interfaces/clk_if.sv"
`include "interfaces/freq_clk_if.sv"
`include "interfaces/i2c_if.sv"
`include "interfaces/irq_if.sv"
`include "interfaces/spi_if.sv"
`include "interfaces/wishbone_if.sv"
`include "interfaces/gmii_if.sv"
`include "interfaces/altera_avalon_mm_if.sv"
`include "interfaces/altera_avalon_st_if.sv"
`include "interfaces/amba_atb_if.sv"
