`include "avlst_uvc/avlst_common.svh"
`include "avlst_uvc/avlst_transaction.svh"
`include "avlst_uvc/avlst_config.svh"
`include "avlst_uvc/avlst_adapter.svh"
`include "avlst_uvc/avlst_sequencer.svh"
`include "avlst_uvc/avlst_driver.svh"
`include "avlst_uvc/avlst_monitor.svh"
`include "avlst_uvc/avlst_agent.svh"
`include "avlst_uvc/avlst_sequence.svh"
