
//------------------------------------------------------------------------------
// Package: test_pkg
//------------------------------------------------------------------------------
package test_pkg;
  `include "uvm_macros.svh"
  import uvm_pkg::*;
  import uvc_pkg::*;
  import toolbox_pkg::*;
  import sknobs::*;
  import tb_pkg::*;
  import sequence_pkg::*;
  
  `include "testcase/base_test.svh"
  `include "testcase/video_file_test.svh"
endpackage : test_pkg
