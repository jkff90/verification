typedef class scb_config;
typedef class scb_txrx_fifo;
typedef class scb_txrx_ooo;
typedef class scb_txrx_ooo_axi;

`include "scb_uvc/scb_common.svh"
`include "scb_uvc/scb_config.svh"
`include "scb_uvc/scb_txrx_fifo.svh"
`include "scb_uvc/scb_txrx_ooo.svh"
`include "scb_uvc/scb_txrx_ooo_axi.svh"
