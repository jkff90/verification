//IP Functional Simulation Model
//VERSION_BEGIN 13.0 cbx_mgl 2013:04:24:18:11:10:SJ cbx_simgen 2013:04:24:18:08:47:SJ  VERSION_END
// synthesis VERILOG_INPUT_VERSION VERILOG_2001
// altera message_off 10463



// Copyright (C) 1991-2013 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.

// You may only use these simulation model output files for simulation
// purposes and expressly not for synthesis or any other purposes (in which
// event Altera disclaims all warranties of any kind).


//synopsys translate_off

//synthesis_resources = altmult_add 6 altsyncram 1 lpm_counter 2 lut 1110 mux21 833 oper_add 30 oper_less_than 1 oper_mux 111 oper_selector 152 
`timescale 1 ps / 1 ps
module  alpha_mixer
	( 
	alpha_in_0_data,
	alpha_in_0_endofpacket,
	alpha_in_0_ready,
	alpha_in_0_startofpacket,
	alpha_in_0_valid,
	alpha_in_1_data,
	alpha_in_1_endofpacket,
	alpha_in_1_ready,
	alpha_in_1_startofpacket,
	alpha_in_1_valid,
	clock,
	control_av_address,
	control_av_chipselect,
	control_av_readdata,
	control_av_write,
	control_av_writedata,
	din_0_data,
	din_0_endofpacket,
	din_0_ready,
	din_0_startofpacket,
	din_0_valid,
	din_1_data,
	din_1_endofpacket,
	din_1_ready,
	din_1_startofpacket,
	din_1_valid,
	dout_data,
	dout_endofpacket,
	dout_ready,
	dout_startofpacket,
	dout_valid,
	reset) /* synthesis synthesis_clearbox=1 */;
	input   [7:0]  alpha_in_0_data;
	input   alpha_in_0_endofpacket;
	output   alpha_in_0_ready;
	input   alpha_in_0_startofpacket;
	input   alpha_in_0_valid;
	input   [7:0]  alpha_in_1_data;
	input   alpha_in_1_endofpacket;
	output   alpha_in_1_ready;
	input   alpha_in_1_startofpacket;
	input   alpha_in_1_valid;
	input   clock;
	input   [5:0]  control_av_address;
	input   control_av_chipselect;
	output   [15:0]  control_av_readdata;
	input   control_av_write;
	input   [15:0]  control_av_writedata;
	input   [23:0]  din_0_data;
	input   din_0_endofpacket;
	output   din_0_ready;
	input   din_0_startofpacket;
	input   din_0_valid;
	input   [23:0]  din_1_data;
	input   din_1_endofpacket;
	output   din_1_ready;
	input   din_1_startofpacket;
	input   din_1_valid;
	output   [23:0]  dout_data;
	output   dout_endofpacket;
	input   dout_ready;
	output   dout_startofpacket;
	output   dout_valid;
	input   reset;

	wire  [17:0]   wire_nl1Oi1O_result;
	wire  [17:0]   wire_nl1OiiO_result;
	wire  [17:0]   wire_nl1OiOO_result;
	wire  [17:0]   wire_nl1Ol0O_result;
	wire  [17:0]   wire_nl1OllO_result;
	wire  [17:0]   wire_nl1OO1O_result;
	wire  [15:0]   wire_niOl0il_q_a;
	wire  [15:0]   wire_niOl0il_q_b;
	reg	ni1i00l63;
	reg	ni1i00l64;
	reg	ni1i00O61;
	reg	ni1i00O62;
	reg	ni1i01i67;
	reg	ni1i01i68;
	reg	ni1i01O65;
	reg	ni1i01O66;
	reg	ni1i0il59;
	reg	ni1i0il60;
	reg	ni1i0iO57;
	reg	ni1i0iO58;
	reg	ni1i0ll55;
	reg	ni1i0ll56;
	reg	ni1i0Oi53;
	reg	ni1i0Oi54;
	reg	ni1i0Ol51;
	reg	ni1i0Ol52;
	reg	ni1i10O79;
	reg	ni1i10O80;
	reg	ni1i1ii77;
	reg	ni1i1ii78;
	reg	ni1i1li75;
	reg	ni1i1li76;
	reg	ni1i1ll73;
	reg	ni1i1ll74;
	reg	ni1i1Oi71;
	reg	ni1i1Oi72;
	reg	ni1i1Ol69;
	reg	ni1i1Ol70;
	reg	ni1ii1i49;
	reg	ni1ii1i50;
	reg	ni1ii1O47;
	reg	ni1ii1O48;
	reg	ni1iill45;
	reg	ni1iill46;
	reg	ni1il0i41;
	reg	ni1il0i42;
	reg	ni1il0l39;
	reg	ni1il0l40;
	reg	ni1il0O37;
	reg	ni1il0O38;
	reg	ni1il1O43;
	reg	ni1il1O44;
	reg	ni1ilii35;
	reg	ni1ilii36;
	reg	ni1ilil33;
	reg	ni1ilil34;
	reg	ni1iliO31;
	reg	ni1iliO32;
	reg	ni1illi29;
	reg	ni1illi30;
	reg	ni1illl27;
	reg	ni1illl28;
	reg	ni1illO25;
	reg	ni1illO26;
	reg	ni1ilOi23;
	reg	ni1ilOi24;
	reg	ni1ilOl21;
	reg	ni1ilOl22;
	reg	ni1ilOO19;
	reg	ni1ilOO20;
	reg	ni1iO0i11;
	reg	ni1iO0i12;
	reg	ni1iO0l10;
	reg	ni1iO0l9;
	reg	ni1iO0O7;
	reg	ni1iO0O8;
	reg	ni1iO1i17;
	reg	ni1iO1i18;
	reg	ni1iO1l15;
	reg	ni1iO1l16;
	reg	ni1iO1O13;
	reg	ni1iO1O14;
	reg	ni1iOii5;
	reg	ni1iOii6;
	reg	ni1iOil3;
	reg	ni1iOil4;
	reg	ni1iOll1;
	reg	ni1iOll2;
	reg	n100i;
	reg	n100l;
	reg	n100O;
	reg	n101i;
	reg	n101l;
	reg	n101O;
	reg	n10ii;
	reg	n10il;
	reg	n10iO;
	reg	n10li;
	reg	n10ll;
	reg	n10lO;
	reg	n10Oi;
	reg	n10Ol;
	reg	n10OO;
	reg	n110i;
	reg	n110l;
	reg	n110O;
	reg	n111i;
	reg	n111l;
	reg	n111O;
	reg	n11ii;
	reg	n11il;
	reg	n11iO;
	reg	n11li;
	reg	n11ll;
	reg	n11lO;
	reg	n11Oi;
	reg	n11Ol;
	reg	n11OO;
	reg	n1i0i;
	reg	n1i0l;
	reg	n1i0O;
	reg	n1i1i;
	reg	n1i1l;
	reg	n1i1O;
	reg	n1iii;
	reg	n1iil;
	reg	n1ili;
	reg	nlO10l;
	reg	nlOOOi;
	reg	nlOOOl;
	reg	nlOOOO;
	reg	ni0101l;
	reg	ni01lil;
	reg	n000i;
	reg	n000l;
	reg	n000O;
	reg	n001i;
	reg	n001l;
	reg	n001O;
	reg	n00ii;
	reg	n00il;
	reg	n00iO;
	reg	n00li;
	reg	n00ll;
	reg	n00lO;
	reg	n00Oi;
	reg	n00Ol;
	reg	n00OO;
	reg	n010i;
	reg	n010l;
	reg	n010O;
	reg	n011O;
	reg	n01ii;
	reg	n01il;
	reg	n01iO;
	reg	n01li;
	reg	n01ll;
	reg	n01lO;
	reg	n01Oi;
	reg	n01Ol;
	reg	n01OO;
	reg	n0i0i;
	reg	n0i0l;
	reg	n0i0O;
	reg	n0i1i;
	reg	n0i1l;
	reg	n0i1O;
	reg	n0iii;
	reg	n0iil;
	reg	n0iiO;
	reg	n0ili;
	reg	n0ill;
	reg	n0ilO;
	reg	n0iOi;
	reg	n0iOl;
	reg	n0iOO;
	reg	n0l0i;
	reg	n0l0l;
	reg	n0l0O;
	reg	n0l1i;
	reg	n0l1l;
	reg	n0l1O;
	reg	n0lii;
	reg	n0lil;
	reg	n0liO;
	reg	n0lli;
	reg	n0lll;
	reg	n0llO;
	reg	n0lOi;
	reg	n0lOl;
	reg	n0lOO;
	reg	n0O0i;
	reg	n0O0l;
	reg	n0O0O;
	reg	n0O1i;
	reg	n0O1l;
	reg	n0O1O;
	reg	n0Oii;
	reg	n0Oil;
	reg	n0OiO;
	reg	n0Oli;
	reg	n0Oll;
	reg	n0OlO;
	reg	n0OOi;
	reg	n0OOl;
	reg	n0OOO;
	reg	n1ill;
	reg	ni10l;
	reg	ni11i;
	reg	ni11l;
	reg	ni11O;
	reg	ni10i_clk_prev;
	wire	wire_ni10i_CLRN;
	wire	wire_ni10i_PRN;
	reg	nii010i;
	reg	nii010l;
	reg	nii010O;
	reg	nii01ii;
	reg	nii01il;
	reg	nii01li;
	reg	nii00li;
	reg	nii0i0i;
	reg	nii0i0l;
	reg	nii0i0O;
	reg	nii0i1i;
	reg	nii0i1l;
	reg	nii0i1O;
	reg	nii0iii;
	reg	nii0iil;
	reg	nii0iiO;
	reg	nii0ili;
	reg	nii0ill;
	reg	nii0ilO;
	reg	nii0iOi;
	reg	nii0iOl;
	reg	nii0iOO;
	reg	nii0l0i;
	reg	nii0l0l;
	reg	nii0l0O;
	reg	nii0l1i;
	reg	nii0l1l;
	reg	nii0l1O;
	reg	nii0lii;
	reg	nii0lil;
	reg	nii0lli;
	reg	ni0O00i;
	reg	ni0O00l;
	reg	ni0O00O;
	reg	ni0O01i;
	reg	ni0O01l;
	reg	ni0O01O;
	reg	ni0O0ii;
	reg	ni0O0il;
	reg	ni0O0iO;
	reg	ni0O0li;
	reg	ni0O0ll;
	reg	ni0O0lO;
	reg	ni0O0Oi;
	reg	ni0O0Ol;
	reg	ni0O0OO;
	reg	ni0O1iO;
	reg	ni0O1li;
	reg	ni0O1ll;
	reg	ni0O1lO;
	reg	ni0O1Oi;
	reg	ni0O1Ol;
	reg	ni0O1OO;
	reg	ni0Oi0l;
	reg	ni0Oi1i;
	reg	ni0Oi1l;
	reg	nii110i;
	reg	nii100i;
	reg	nii100l;
	reg	nii100O;
	reg	nii101i;
	reg	nii101l;
	reg	nii101O;
	reg	nii10ii;
	reg	nii10il;
	reg	nii10iO;
	reg	nii10li;
	reg	nii10ll;
	reg	nii10lO;
	reg	nii10Oi;
	reg	nii10Ol;
	reg	nii10OO;
	reg	nii11lO;
	reg	nii11Oi;
	reg	nii11Ol;
	reg	nii11OO;
	reg	nii1i0i;
	reg	nii1i0l;
	reg	nii1i1i;
	reg	nii1i1l;
	reg	nii1i1O;
	reg	nii1iii;
	reg	nii1iiO;
	reg	nii1ili;
	reg	nii1ill;
	reg	nii1ilO;
	reg	nii1iOi;
	reg	nii1iOl;
	reg	nii1iOO;
	reg	nii1l0i;
	reg	nii1l1i;
	reg	nii1l1l;
	reg	nii1lii;
	reg	nii1lil;
	reg	nii1liO;
	reg	nii1lli;
	reg	nii1lll;
	reg	nii1llO;
	reg	nii1lOi;
	reg	nii1lOO;
	reg	nii1O0i;
	wire	wire_nii1O1O_ENA;
	reg	nii1Oil;
	reg	nii1OiO;
	reg	nii1Oli;
	reg	nii1OlO;
	reg	nil10lO;
	reg	nil1i0i;
	reg	nil1i0l;
	reg	nil1i0O;
	reg	nil1i1O;
	reg	nil1iii;
	reg	nil1iil;
	reg	nil1iiO;
	reg	nil1ili;
	reg	nil1ill;
	reg	nil1ilO;
	reg	nil1iOi;
	reg	nil1iOl;
	reg	nil1iOO;
	reg	nil1l0i;
	reg	nil1l0l;
	reg	nil1l0O;
	reg	nil1l1i;
	reg	nil1l1l;
	reg	nil1l1O;
	reg	nil1lii;
	reg	nil1lil;
	reg	nil1liO;
	reg	nil1lli;
	reg	nil1llO;
	reg	nilOiOl;
	reg	nilOl0l;
	reg	nilOl0O;
	reg	nilOlii;
	reg	nilOlil;
	reg	nilOliO;
	reg	nilOlli;
	reg	nilOlll;
	reg	nilOlOi;
	reg	niOii1l;
	wire	wire_niOii1i_ENA;
	reg	niOii0i;
	reg	niOiill;
	reg	niOiilO;
	reg	niOiiOi;
	reg	niOiiOl;
	reg	niOiiOO;
	reg	niOil0i;
	reg	niOil0l;
	reg	niOil0O;
	reg	niOil1i;
	reg	niOil1l;
	reg	niOil1O;
	reg	niOilii;
	reg	niOilil;
	reg	niOiliO;
	reg	niOilli;
	reg	niOilll;
	reg	niOillO;
	reg	niOilOi;
	reg	niOilOl;
	reg	niOilOO;
	reg	niOiO0l;
	reg	niOiO1i;
	reg	niOiO1l;
	reg	niOiO1O;
	reg	ni0000l;
	reg	ni0001i;
	reg	ni0001O;
	reg	ni000il;
	reg	ni000li;
	reg	ni000lO;
	reg	ni0011l;
	reg	ni001ii;
	reg	ni001ll;
	reg	ni001Ol;
	reg	ni00i0O;
	reg	ni00i1l;
	reg	ni00iiO;
	reg	ni00ill;
	reg	ni00iOi;
	reg	ni00iOO;
	reg	ni00l0l;
	reg	ni00l1O;
	reg	ni00lii;
	reg	ni00llO;
	reg	ni00O0i;
	reg	ni00O0O;
	reg	ni00O1i;
	reg	ni00Oil;
	reg	ni0100l;
	reg	ni010ii;
	reg	ni01i1O;
	reg	ni01iii;
	reg	ni01iil;
	reg	ni01liO;
	reg	ni01lli;
	reg	ni01Oli;
	reg	ni01OOi;
	reg	ni01OOO;
	reg	ni0Oi0i;
	reg	ni0Oi1O;
	reg	nii0lll;
	reg	nii0lOi;
	reg	nii0lOl;
	reg	nii0lOO;
	reg	nii0O0i;
	reg	nii0O0l;
	reg	nii0O0O;
	reg	nii0O1i;
	reg	nii0O1l;
	reg	nii0O1O;
	reg	nii0Oii;
	reg	nii0Oil;
	reg	nii0OiO;
	reg	nii0Oli;
	reg	nii0Oll;
	reg	nii0OlO;
	reg	nii0OOi;
	reg	nii0OOl;
	reg	nii0OOO;
	reg	niii00i;
	reg	niii00l;
	reg	niii00O;
	reg	niii01i;
	reg	niii01l;
	reg	niii01O;
	reg	niii0ii;
	reg	niii0il;
	reg	niii0iO;
	reg	niii0li;
	reg	niii0ll;
	reg	niii0lO;
	reg	niii0Oi;
	reg	niii0Ol;
	reg	niii0OO;
	reg	niii10i;
	reg	niii10l;
	reg	niii10O;
	reg	niii11i;
	reg	niii11l;
	reg	niii11O;
	reg	niii1ii;
	reg	niii1il;
	reg	niii1iO;
	reg	niii1li;
	reg	niii1ll;
	reg	niii1lO;
	reg	niii1Oi;
	reg	niii1Ol;
	reg	niii1OO;
	reg	niiii0i;
	reg	niiii0l;
	reg	niiii0O;
	reg	niiii1i;
	reg	niiii1l;
	reg	niiii1O;
	reg	niiiiii;
	reg	niiiiil;
	reg	niiiiiO;
	reg	niiiili;
	reg	niiiill;
	reg	niiiilO;
	reg	niiiiOi;
	reg	niiiiOl;
	reg	niiiiOO;
	reg	niiil0i;
	reg	niiil0l;
	reg	niiil0O;
	reg	niiil1i;
	reg	niiil1l;
	reg	niiil1O;
	reg	niiilii;
	reg	niiilil;
	reg	niiiliO;
	reg	niiilli;
	reg	niiilll;
	reg	niiillO;
	reg	niiilOi;
	reg	niiilOl;
	reg	nil000i;
	reg	nil000l;
	reg	nil000O;
	reg	nil001i;
	reg	nil001l;
	reg	nil001O;
	reg	nil00ii;
	reg	nil00il;
	reg	nil00iO;
	reg	nil00li;
	reg	nil00ll;
	reg	nil00lO;
	reg	nil00Oi;
	reg	nil00Ol;
	reg	nil00OO;
	reg	nil010i;
	reg	nil010l;
	reg	nil010O;
	reg	nil011i;
	reg	nil011l;
	reg	nil011O;
	reg	nil01ii;
	reg	nil01il;
	reg	nil01iO;
	reg	nil01li;
	reg	nil01ll;
	reg	nil01lO;
	reg	nil01Oi;
	reg	nil01Ol;
	reg	nil01OO;
	reg	nil0i0i;
	reg	nil0i0l;
	reg	nil0i0O;
	reg	nil0i1i;
	reg	nil0i1l;
	reg	nil0i1O;
	reg	nil0iii;
	reg	nil0iil;
	reg	nil0iiO;
	reg	nil0ili;
	reg	nil0ill;
	reg	nil0ilO;
	reg	nil0iOi;
	reg	nil0iOl;
	reg	nil0iOO;
	reg	nil0l0i;
	reg	nil0l0l;
	reg	nil0l0O;
	reg	nil0l1i;
	reg	nil0l1l;
	reg	nil0l1O;
	reg	nil0lii;
	reg	nil0lil;
	reg	nil0liO;
	reg	nil0lli;
	reg	nil0lll;
	reg	nil0llO;
	reg	nil0lOi;
	reg	nil0lOl;
	reg	nil0lOO;
	reg	nil0O1i;
	reg	nil101O;
	reg	nil11Ol;
	reg	nil11OO;
	reg	nil1lOi;
	reg	nil1lOO;
	reg	nil1O0i;
	reg	nil1O0l;
	reg	nil1O0O;
	reg	nil1O1i;
	reg	nil1O1l;
	reg	nil1O1O;
	reg	nil1Oii;
	reg	nil1Oil;
	reg	nil1OiO;
	reg	nil1Oli;
	reg	nil1Oll;
	reg	nil1OlO;
	reg	nil1OOi;
	reg	nil1OOl;
	reg	nil1OOO;
	reg	nilO00l;
	reg	nilO01i;
	reg	nilO01l;
	reg	nilO0iO;
	reg	nilO0li;
	reg	nilO0ll;
	reg	nilOi0l;
	reg	nilOlOl;
	reg	nilOO0i;
	reg	nilOO0l;
	reg	nilOO0O;
	reg	nilOO1i;
	reg	nilOO1l;
	reg	nilOO1O;
	reg	nilOOii;
	reg	nilOOil;
	reg	nilOOiO;
	reg	nilOOli;
	reg	nilOOll;
	reg	nilOOlO;
	reg	nilOOOi;
	reg	nilOOOl;
	reg	nilOOOO;
	reg	niO00il;
	reg	niO00iO;
	reg	niO00lO;
	reg	niO110i;
	reg	niO110l;
	reg	niO110O;
	reg	niO111i;
	reg	niO111l;
	reg	niO111O;
	reg	niO11ii;
	reg	niO11il;
	reg	niO11iO;
	reg	niO11li;
	reg	niO11ll;
	reg	niO11lO;
	reg	niO11Oi;
	reg	niO11Ol;
	reg	niOii0l;
	reg	niOiOii;
	reg	niOl0Ol;
	reg	niOl0OO;
	reg	niOli0i;
	reg	niOli0l;
	reg	niOli0O;
	reg	niOli1i;
	reg	niOli1l;
	reg	niOli1O;
	reg	niOliii;
	reg	niOliil;
	reg	niOlili;
	reg	niOlO0i;
	reg	niOlO0l;
	reg	niOlO0O;
	reg	niOlO1l;
	reg	niOlO1O;
	reg	niOlOii;
	reg	niOlOil;
	reg	niOlOiO;
	reg	niOlOli;
	reg	niOlOlO;
	reg	niOO00i;
	reg	niOO00l;
	reg	niOO01i;
	reg	niOO01l;
	reg	niOO01O;
	reg	niOO0ii;
	reg	niOO1Ol;
	reg	niOO1OO;
	reg	niOO10i;
	reg	niOO10l;
	reg	niOO10O;
	reg	niOO11i;
	reg	niOO11l;
	reg	niOO11O;
	reg	niOO1ii;
	reg	niOO1il;
	reg	niOO1iO;
	reg	niOO1ll;
	reg	niOO0ll;
	reg	niOO0lO;
	reg	niOO0Oi;
	reg	niOO0Ol;
	reg	niOO0OO;
	reg	niOOi0i;
	reg	niOOi1i;
	reg	niOOi1l;
	reg	nl00i0l;
	reg	nl00i0O;
	reg	nl00iii;
	reg	nl00iil;
	reg	nl00iiO;
	reg	nl00ili;
	reg	nl00ill;
	reg	nl00ilO;
	reg	nl00iOi;
	reg	nl00iOO;
	reg	nl00l0i;
	reg	nl00l0l;
	reg	nl00l0O;
	reg	nl00l1l;
	reg	nl00l1O;
	reg	nl00lil;
	reg	nl00lli;
	wire	wire_nl00liO_ENA;
	reg	nl00llO;
	reg	nl00lOi;
	reg	nl00lOl;
	reg	nl00O1i;
	reg	nl00O0i;
	wire	wire_nl00O1O_ENA;
	reg	nl00O0O;
	reg	nl00Oii;
	reg	nl00Oil;
	reg	nl00Oli;
	reg	nl0100i;
	reg	nl0100O;
	reg	nl0101l;
	reg	nl0101O;
	reg	nl0110l;
	reg	nl011ii;
	reg	nl01i0l;
	reg	nl01i1i;
	reg	nl01i1l;
	reg	nl01i1O;
	reg	nl0i0ll;
	reg	nl0i0Oi;
	wire	wire_nl0i0lO_ENA;
	reg	nl0i10l;
	reg	nl00OlO;
	reg	nl00OOi;
	reg	nl00OOl;
	reg	nl00OOO;
	reg	nl0i11i;
	reg	nl0i11O;
	reg	nl0i10O;
	reg	nl0i1ii;
	reg	nl0i1il;
	reg	nl0i1iO;
	reg	nl0i1li;
	reg	nl0i1ll;
	reg	nl0i1lO;
	reg	nl0i1Ol;
	reg	nl0i0OO;
	reg	nl0ii0i;
	reg	nl0ii0l;
	reg	nl0ii0O;
	reg	nl0ii1i;
	reg	nl0ii1l;
	reg	nl0ii1O;
	reg	nl0iiii;
	reg	nl0iiil;
	reg	nl0iili;
	reg	nl0ilil;
	reg	nl0iliO;
	reg	nl0illi;
	reg	nl0illl;
	reg	nl0illO;
	reg	nl0ilOi;
	reg	nl0ilOl;
	reg	nl0ilOO;
	reg	nl0iO1i;
	reg	nl0iO1O;
	reg	nl0l0il;
	wire	wire_nl0l0ii_ENA;
	reg	nl0l0Oi;
	wire	wire_nl0l0lO_ENA;
	reg	nl0li1i;
	wire	wire_nl0l0OO_ENA;
	reg	nl0l10l;
	wire	wire_nl0l10i_ENA;
	reg	nl0l11l;
	wire	wire_nl0l11i_ENA;
	reg	nl0l1il;
	wire	wire_nl0l1ii_ENA;
	reg	nl0l1ll;
	wire	wire_nl0l1li_ENA;
	reg	nl0l1Oi;
	reg	nl0l1OO;
	reg	nl0liii;
	wire	wire_nl0li0O_ENA;
	reg	nl0li0i;
	wire	wire_nl0li1O_ENA;
	reg	nl0lili;
	wire	wire_nl0liiO_ENA;
	reg	nl0lO0i;
	reg	nl0lO0l;
	reg	nl0lO0O;
	reg	nl0lOii;
	reg	nl0lOil;
	reg	nl0lOiO;
	reg	nl0lOli;
	reg	nl0lOll;
	reg	nl0lOlO;
	reg	nl0lOOi;
	reg	nl0lOOO;
	reg	nl0O01i;
	wire	wire_nl0O1OO_ENA;
	reg	nl0OiOl;
	reg	nl0OiOO;
	reg	nl0Ol0i;
	reg	nl0Ol0l;
	reg	nl0Ol1i;
	reg	nl0Ol1l;
	reg	nl0Ol1O;
	reg	nl0Olii;
	reg	nl100iO;
	reg	nl100li;
	reg	nl100ll;
	reg	nl100lO;
	reg	nl100Oi;
	reg	nl100Ol;
	reg	nl100OO;
	reg	nl10i0i;
	reg	nl10i0l;
	reg	nl10i0O;
	reg	nl10i1i;
	reg	nl10i1l;
	reg	nl10i1O;
	reg	nl10iii;
	reg	nl10iil;
	reg	nl10iiO;
	reg	nl10ili;
	reg	nl10ill;
	reg	nl10ilO;
	reg	nl10iOi;
	reg	nl10iOl;
	reg	nl10iOO;
	reg	nl10l1i;
	reg	nl10l1O;
	reg	nl10llO;
	reg	nl10lOO;
	reg	nl10l0O;
	reg	nl10lii;
	reg	nl10lil;
	reg	nl10liO;
	reg	nl10lli;
	reg	nl10lll;
	reg	nl10lOi;
	reg	nl10O1l;
	reg	nl10Oll;
	reg	nl10OOl;
	reg	nl10O0l;
	reg	nl10O0O;
	reg	nl10Oii;
	reg	nl10Oil;
	reg	nl10OiO;
	reg	nl10Oli;
	reg	nl10OlO;
	reg	nl1i11i;
	reg	nl1100i;
	reg	nl1100l;
	reg	nl1100O;
	reg	nl1101l;
	reg	nl1101O;
	reg	nl110ii;
	reg	nl110il;
	reg	nl110iO;
	reg	nl110li;
	reg	nl110ll;
	reg	nl110lO;
	reg	nl110Oi;
	reg	nl110Ol;
	reg	nl110OO;
	reg	nl11i0i;
	reg	nl11i0l;
	reg	nl11i0O;
	reg	nl11i1i;
	reg	nl11i1l;
	reg	nl11i1O;
	reg	nl11iii;
	reg	nl11iil;
	reg	nl11iiO;
	reg	nl11ill;
	reg	nl1i00l;
	reg	nl1i01i;
	reg	nl1i01l;
	reg	nl1i01O;
	reg	nl1i00O;
	reg	nl1i0ii;
	reg	nl1i0il;
	reg	nl1i0li;
	reg	nl1i0Oi;
	reg	nl1i0OO;
	reg	nl1i10i;
	reg	nl1i10l;
	reg	nl1i10O;
	reg	nl1i1il;
	reg	nl1i1iO;
	reg	nl1i1li;
	reg	nl1i1ll;
	reg	nl1i1Oi;
	reg	nl1ii0i;
	reg	nl1ii0l;
	reg	nl1ii0O;
	reg	nl1ii1l;
	reg	nl1ii1O;
	reg	nl1iiii;
	reg	nl1iiil;
	reg	nl1iili;
	reg	nl1iilO;
	reg	nl1iiOi;
	reg	nl1iiOl;
	reg	nl1iiOO;
	reg	nl1il0l;
	reg	nl1il1i;
	reg	nl1il1l;
	reg	nl1il1O;
	reg	nl1ilii;
	reg	nl1ilil;
	reg	nl1iliO;
	reg	nl1illi;
	reg	nl1illl;
	reg	nl1illO;
	reg	nl1ilOi;
	reg	nl1ilOO;
	reg	nl1iO0i;
	reg	nl1iO0l;
	reg	nl1iO0O;
	reg	nl1iO1l;
	reg	nl1iO1O;
	reg	nl1iOii;
	reg	nl1iOil;
	reg	nl1iOli;
	reg	nl1l01l;
	reg	nl1l1iO;
	reg	nl1l1li;
	reg	nl1l1ll;
	reg	nl1l1lO;
	reg	nl1l1Oi;
	reg	nl1l1Ol;
	reg	nl1l1OO;
	reg	nl1iOOi;
	reg	nl1iOOl;
	reg	nl1iOOO;
	reg	nl1l10i;
	reg	nl1l10O;
	reg	nl1l11i;
	reg	nl1l11l;
	reg	nl1l11O;
	reg	nl1llll;
	reg	nl1lllO;
	reg	nl1llOi;
	reg	nl1llOl;
	reg	nl1llOO;
	reg	nl1lO0i;
	reg	nl1lO1i;
	reg	nl1lO1l;
	reg	nl1O00i;
	reg	nl1O00O;
	reg	nl1O01i;
	reg	nl1O01l;
	reg	nl1O01O;
	reg	nl1O1lO;
	reg	nl1O1Oi;
	reg	nl1O1Ol;
	reg	nl1O1OO;
	reg	nl1O10i;
	reg	nl1O10l;
	reg	nl1O10O;
	reg	nl1O11i;
	reg	nl1O11l;
	reg	nl1O11O;
	reg	nl1O1ii;
	reg	nl1O1il;
	reg	nl1O1li;
	reg	niiilOO;
	reg	nil0O1l;
	reg	niO11OO;
	reg	nl1Oi0i;
	reg	nl1Oiil;
	reg	nl1Oili;
	reg	nl1OiOl;
	reg	nl1Ol0l;
	reg	nl1Ol1i;
	reg	nl1Olii;
	reg	nl1Olll;
	reg	nl1OlOi;
	reg	nl1OO0i;
	reg	nl1OO1l;
	reg	nl1OOiO;
	reg	nl1OOll;
	wire	wire_nl1OOli_ENA;
	reg	nl1OOOl;
	wire	wire_nl1OOOi_ENA;
	reg	nli000l;
	reg	nli001i;
	reg	nli001l;
	reg	nli001O;
	reg	nli01lO;
	reg	nli01Oi;
	reg	nli01Ol;
	reg	nli01OO;
	wire	wire_nli000i_CLRN;
	reg	nli00ii;
	reg	nli00il;
	reg	nli00iO;
	reg	nli00li;
	reg	nli00ll;
	reg	nli00lO;
	reg	nli00Oi;
	reg	nli00OO;
	reg	nli00Ol_clk_prev;
	wire	wire_nli00Ol_CLRN;
	wire	wire_nli00Ol_PRN;
	reg	nli010i;
	reg	nli010l;
	reg	nli010O;
	reg	nli011l;
	reg	nli011O;
	reg	nli01ii;
	reg	nli01il;
	reg	nli01li;
	reg	nli01iO_clk_prev;
	wire	wire_nli01iO_PRN;
	reg	nli0i0i;
	reg	nli0i0l;
	reg	nli0i0O;
	reg	nli0i1l;
	reg	nli0i1O;
	reg	nli0iii;
	reg	nli0iil;
	reg	nli0ili;
	reg	nli0iiO_clk_prev;
	wire	wire_nli0iiO_CLRN;
	wire	wire_nli0iiO_PRN;
	reg	nli0ilO;
	reg	nli0iOi;
	reg	nli0iOl;
	reg	nli0iOO;
	reg	nli0l0l;
	reg	nli0l1i;
	reg	nli0l1l;
	reg	nli0l1O;
	wire	wire_nli0l0i_CLRN;
	reg	nli0lii;
	reg	nli0lil;
	reg	nli0liO;
	reg	nli0lli;
	reg	nli0lll;
	reg	nli0llO;
	reg	nli0lOi;
	reg	nli0lOO;
	reg	nli0lOl_clk_prev;
	wire	wire_nli0lOl_CLRN;
	wire	wire_nli0lOl_PRN;
	reg	nli100O;
	wire	wire_nli100l_ENA;
	reg	nli101O;
	wire	wire_nli101l_ENA;
	reg	nli10iO;
	wire	wire_nli10il_ENA;
	reg	nli10lO;
	wire	wire_nli10ll_ENA;
	reg	nli10OO;
	wire	wire_nli10Ol_ENA;
	reg	nli11lO;
	wire	wire_nli11ll_ENA;
	reg	nli11OO;
	wire	wire_nli11Ol_ENA;
	reg	nli1i0O;
	wire	wire_nli1i0l_ENA;
	reg	nli1i1O;
	wire	wire_nli1i1l_ENA;
	reg	nli1iiO;
	wire	wire_nli1iil_ENA;
	reg	nli1ilO;
	wire	wire_nli1ill_CLRN;
	wire	wire_nli1ill_ENA;
	reg	nli1iOO;
	wire	wire_nli1iOl_CLRN;
	wire	wire_nli1iOl_ENA;
	reg	nli1l0i;
	reg	nli1l0l;
	reg	nli1l0O;
	reg	nli1l1l;
	reg	nli1l1O;
	reg	nli1lii;
	reg	nli1lil;
	reg	nli1lli;
	reg	nli1llO;
	reg	nli1lOi;
	reg	nli1lOl;
	reg	nli1lOO;
	reg	nli1O0l;
	reg	nli1O1i;
	reg	nli1O1l;
	reg	nli1O1O;
	reg	nli1O0i_clk_prev;
	wire	wire_nli1O0i_CLRN;
	wire	wire_nli1O0i_PRN;
	reg	nli1Oii;
	reg	nli1Oil;
	reg	nli1OiO;
	reg	nli1Oli;
	reg	nli1Oll;
	reg	nli1OlO;
	reg	nli1OOi;
	reg	nli1OOO;
	reg	nli1OOl_clk_prev;
	wire	wire_nli1OOl_CLRN;
	wire	wire_nli1OOl_PRN;
	reg	nlii00l;
	reg	nlii01i;
	reg	nlii01l;
	reg	nlii01O;
	wire	wire_nlii00i_CLRN;
	reg	nlii0ii;
	reg	nlii0il;
	reg	nlii0iO;
	reg	nlii0ll;
	reg	nli0O0i;
	reg	nli0O0l;
	reg	nli0O0O;
	reg	nli0O1l;
	reg	nli0O1O;
	reg	nli0Oii;
	reg	nli0Oil;
	reg	nli0OiO;
	reg	nli0Oli;
	reg	nli0Oll;
	reg	nli0OlO;
	reg	nli0OOi;
	reg	nli0OOl;
	reg	nli0OOO;
	reg	nlii10i;
	reg	nlii10l;
	reg	nlii10O;
	reg	nlii11i;
	reg	nlii11l;
	reg	nlii11O;
	reg	nlii1ii;
	reg	nlii1il;
	reg	nlii1iO;
	reg	nlii1ll;
	reg	nlii1li_clk_prev;
	wire	wire_nlii1li_PRN;
	reg	nlii1Ol;
	wire	wire_nlii1Oi_ENA;
	reg	nlii0Oi;
	reg	nlii0Ol;
	reg	nlii0OO;
	reg	nliii1l;
	reg	ni0000i;
	reg	ni0000O;
	reg	ni0001l;
	reg	ni000ii;
	reg	ni000iO;
	reg	ni000ll;
	reg	ni000Oi;
	reg	ni000Ol;
	reg	ni000OO;
	reg	ni0010i;
	reg	ni0010l;
	reg	ni0010O;
	reg	ni0011i;
	reg	ni0011O;
	reg	ni001il;
	reg	ni001iO;
	reg	ni001li;
	reg	ni001lO;
	reg	ni001Oi;
	reg	ni001OO;
	reg	ni00i0i;
	reg	ni00i0l;
	reg	ni00i1i;
	reg	ni00i1O;
	reg	ni00iii;
	reg	ni00iil;
	reg	ni00ili;
	reg	ni00ilO;
	reg	ni00iOl;
	reg	ni00l0i;
	reg	ni00l0O;
	reg	ni00l1i;
	reg	ni00l1l;
	reg	ni00lil;
	reg	ni00liO;
	reg	ni00lli;
	reg	ni00lll;
	reg	ni00lOi;
	reg	ni00lOl;
	reg	ni00lOO;
	reg	ni00O0l;
	reg	ni00O1l;
	reg	ni00O1O;
	reg	ni00Oii;
	reg	ni0100O;
	reg	ni01Oll;
	reg	ni01OlO;
	reg	ni01OOl;
	reg	ni0il1O;
	reg	nl001li;
	reg	nl001ll;
	reg	nl01O0l;
	reg	nl01O0O;
	reg	nllOOO;
	reg	nlO1Oi;
	reg	nlO1lO_clk_prev;
	wire	wire_nlO1lO_CLRN;
	wire  [6:0]   wire_nl001iO_q;
	wire  [7:0]   wire_nl01O0i_q;
	wire	wire_ni00OiO_dataout;
	wire	wire_ni00Oli_dataout;
	wire	wire_ni00Oll_dataout;
	wire	wire_ni00OlO_dataout;
	wire	wire_ni00OOi_dataout;
	wire	wire_ni00OOl_dataout;
	wire	wire_ni00OOO_dataout;
	wire	wire_ni010il_dataout;
	wire	wire_ni010iO_dataout;
	wire	wire_ni010li_dataout;
	wire	wire_ni010ll_dataout;
	wire	wire_ni010lO_dataout;
	wire	wire_ni010Oi_dataout;
	wire	wire_ni0111i_dataout;
	wire	wire_ni0111l_dataout;
	wire	wire_ni01i0i_dataout;
	wire	wire_ni01iiO_dataout;
	wire	wire_ni01ili_dataout;
	wire	wire_ni01ill_dataout;
	wire	wire_ni01ilO_dataout;
	wire	wire_ni01iOi_dataout;
	wire	wire_ni01iOl_dataout;
	wire	wire_ni01l1i_dataout;
	wire	wire_ni01lll_dataout;
	wire	wire_ni01llO_dataout;
	wire	wire_ni01lOi_dataout;
	wire	wire_ni01lOl_dataout;
	wire	wire_ni0i00i_dataout;
	wire	wire_ni0i00l_dataout;
	wire	wire_ni0i00O_dataout;
	wire	wire_ni0i01i_dataout;
	wire	wire_ni0i01l_dataout;
	wire	wire_ni0i01O_dataout;
	wire	wire_ni0i0ii_dataout;
	wire	wire_ni0i0il_dataout;
	wire	wire_ni0i0iO_dataout;
	wire	wire_ni0i0li_dataout;
	wire	wire_ni0i0ll_dataout;
	wire	wire_ni0i0lO_dataout;
	wire	wire_ni0i0Oi_dataout;
	wire	wire_ni0i0Ol_dataout;
	wire	wire_ni0i0OO_dataout;
	wire	wire_ni0i10i_dataout;
	wire	wire_ni0i10l_dataout;
	wire	wire_ni0i10O_dataout;
	wire	wire_ni0i11i_dataout;
	wire	wire_ni0i11l_dataout;
	wire	wire_ni0i11O_dataout;
	wire	wire_ni0i1ii_dataout;
	wire	wire_ni0i1il_dataout;
	wire	wire_ni0i1iO_dataout;
	wire	wire_ni0i1li_dataout;
	wire	wire_ni0i1ll_dataout;
	wire	wire_ni0i1lO_dataout;
	wire	wire_ni0i1Oi_dataout;
	wire	wire_ni0i1Ol_dataout;
	wire	wire_ni0i1OO_dataout;
	wire	wire_ni0ii0i_dataout;
	wire	wire_ni0ii0l_dataout;
	wire	wire_ni0ii0O_dataout;
	wire	wire_ni0ii1i_dataout;
	wire	wire_ni0ii1l_dataout;
	wire	wire_ni0ii1O_dataout;
	wire	wire_ni0iiii_dataout;
	wire	wire_ni0iiil_dataout;
	wire	wire_ni0iiiO_dataout;
	wire	wire_ni0iili_dataout;
	wire	wire_ni0iill_dataout;
	wire	wire_ni0iilO_dataout;
	wire	wire_ni0iiOi_dataout;
	wire	wire_ni0il0i_dataout;
	wire	wire_ni0il0l_dataout;
	wire	wire_ni0il0O_dataout;
	wire	wire_ni0ilii_dataout;
	wire	wire_ni0ilil_dataout;
	wire	wire_ni0iliO_dataout;
	wire	wire_ni0illi_dataout;
	wire	wire_ni0illl_dataout;
	wire	wire_ni0illO_dataout;
	wire	wire_ni0ilOi_dataout;
	wire	wire_ni0ilOl_dataout;
	wire	wire_ni0ilOO_dataout;
	wire	wire_ni0iO0i_dataout;
	wire	wire_ni0iO0l_dataout;
	wire	wire_ni0iO0O_dataout;
	wire	wire_ni0iO1i_dataout;
	wire	wire_ni0iO1l_dataout;
	wire	wire_ni0iO1O_dataout;
	wire	wire_ni0iOii_dataout;
	wire	wire_ni0iOil_dataout;
	wire	wire_ni0iOiO_dataout;
	wire	wire_ni0iOli_dataout;
	wire	wire_ni0iOll_dataout;
	wire	wire_ni0iOlO_dataout;
	wire	wire_ni0iOOi_dataout;
	wire	wire_ni0iOOl_dataout;
	wire	wire_ni0iOOO_dataout;
	wire	wire_ni0l00i_dataout;
	wire	wire_ni0l00l_dataout;
	wire	wire_ni0l00O_dataout;
	wire	wire_ni0l01i_dataout;
	wire	wire_ni0l01l_dataout;
	wire	wire_ni0l01O_dataout;
	wire	wire_ni0l0ii_dataout;
	wire	wire_ni0l0il_dataout;
	wire	wire_ni0l0Oi_dataout;
	wire	wire_ni0l0Ol_dataout;
	wire	wire_ni0l0OO_dataout;
	wire	wire_ni0l10i_dataout;
	wire	wire_ni0l10l_dataout;
	wire	wire_ni0l10O_dataout;
	wire	wire_ni0l11i_dataout;
	wire	wire_ni0l11l_dataout;
	wire	wire_ni0l11O_dataout;
	wire	wire_ni0l1ii_dataout;
	wire	wire_ni0l1il_dataout;
	wire	wire_ni0l1iO_dataout;
	wire	wire_ni0l1li_dataout;
	wire	wire_ni0l1ll_dataout;
	wire	wire_ni0l1lO_dataout;
	wire	wire_ni0l1Oi_dataout;
	wire	wire_ni0l1Ol_dataout;
	wire	wire_ni0l1OO_dataout;
	wire	wire_ni0li0i_dataout;
	wire	wire_ni0li0l_dataout;
	wire	wire_ni0li0O_dataout;
	wire	wire_ni0li1i_dataout;
	wire	wire_ni0li1l_dataout;
	wire	wire_ni0li1O_dataout;
	wire	wire_ni0liii_dataout;
	wire	wire_ni0liil_dataout;
	wire	wire_ni0liiO_dataout;
	wire	wire_ni0lili_dataout;
	wire	wire_ni0lill_dataout;
	wire	wire_ni0lilO_dataout;
	wire	wire_ni0liOi_dataout;
	wire	wire_ni0liOl_dataout;
	wire	wire_ni0liOO_dataout;
	wire	wire_ni0ll0i_dataout;
	wire	wire_ni0ll0l_dataout;
	wire	wire_ni0ll0O_dataout;
	wire	wire_ni0ll1i_dataout;
	wire	wire_ni0ll1l_dataout;
	wire	wire_ni0ll1O_dataout;
	wire	wire_ni0llii_dataout;
	wire	wire_ni0llil_dataout;
	wire	wire_ni0lliO_dataout;
	wire	wire_ni0llli_dataout;
	wire	wire_ni0llll_dataout;
	wire	wire_ni0lllO_dataout;
	wire	wire_ni0llOi_dataout;
	wire	wire_ni0llOl_dataout;
	wire	wire_ni0llOO_dataout;
	wire	wire_ni0lO0i_dataout;
	wire	wire_ni0lO0l_dataout;
	wire	wire_ni0lO0O_dataout;
	wire	wire_ni0lO1i_dataout;
	wire	wire_ni0lO1l_dataout;
	wire	wire_ni0lO1O_dataout;
	wire	wire_ni0lOii_dataout;
	wire	wire_ni0lOil_dataout;
	wire	wire_ni0lOiO_dataout;
	wire	wire_ni0lOli_dataout;
	wire	wire_ni0lOll_dataout;
	wire	wire_ni0lOlO_dataout;
	wire	wire_ni0lOOi_dataout;
	wire	wire_ni0lOOl_dataout;
	wire	wire_ni0lOOO_dataout;
	wire	wire_ni0O11i_dataout;
	wire	wire_ni0O11l_dataout;
	wire	wire_ni0O1il_dataout;
	wire	wire_ni0Oi0O_dataout;
	wire	wire_ni0Oiii_dataout;
	wire	wire_ni0OilO_dataout;
	wire	wire_ni0OiOi_dataout;
	wire	wire_ni0OiOl_dataout;
	wire	wire_ni0OiOO_dataout;
	wire	wire_ni0Ol0i_dataout;
	wire	wire_ni0Ol0l_dataout;
	wire	wire_ni0Ol0O_dataout;
	wire	wire_ni0Ol1i_dataout;
	wire	wire_ni0Ol1l_dataout;
	wire	wire_ni0Ol1O_dataout;
	wire	wire_ni0Olii_dataout;
	wire	wire_ni0Olil_dataout;
	wire	wire_ni0OliO_dataout;
	wire	wire_ni0Olli_dataout;
	wire	wire_ni0Olll_dataout;
	wire	wire_ni0OllO_dataout;
	wire	wire_ni0OlOi_dataout;
	wire	wire_ni0OlOl_dataout;
	wire	wire_ni0OlOO_dataout;
	wire	wire_ni0OO0i_dataout;
	wire	wire_ni0OO0l_dataout;
	wire	wire_ni0OO0O_dataout;
	wire	wire_ni0OO1i_dataout;
	wire	wire_ni0OO1l_dataout;
	wire	wire_ni0OO1O_dataout;
	wire	wire_ni1l00i_dataout;
	wire	wire_ni1l00l_dataout;
	wire	wire_ni1l00O_dataout;
	wire	wire_ni1l01i_dataout;
	wire	wire_ni1l01l_dataout;
	wire	wire_ni1l01O_dataout;
	wire	wire_ni1l0ii_dataout;
	wire	wire_ni1l0il_dataout;
	wire	wire_ni1l0iO_dataout;
	wire	wire_ni1l0li_dataout;
	wire	wire_ni1l0ll_dataout;
	wire	wire_ni1l0lO_dataout;
	wire	wire_ni1l0Oi_dataout;
	wire	wire_ni1l0Ol_dataout;
	wire	wire_ni1l0OO_dataout;
	wire	wire_ni1l10i_dataout;
	wire	wire_ni1l10l_dataout;
	wire	wire_ni1l10O_dataout;
	wire	wire_ni1l11O_dataout;
	wire	wire_ni1l1ii_dataout;
	wire	wire_ni1l1il_dataout;
	wire	wire_ni1l1iO_dataout;
	wire	wire_ni1l1li_dataout;
	wire	wire_ni1l1ll_dataout;
	wire	wire_ni1l1lO_dataout;
	wire	wire_ni1l1Oi_dataout;
	wire	wire_ni1l1Ol_dataout;
	wire	wire_ni1l1OO_dataout;
	wire	wire_ni1li0i_dataout;
	wire	wire_ni1li0l_dataout;
	wire	wire_ni1li0O_dataout;
	wire	wire_ni1li1i_dataout;
	wire	wire_ni1li1l_dataout;
	wire	wire_ni1li1O_dataout;
	wire	wire_ni1liii_dataout;
	wire	wire_ni1liil_dataout;
	wire	wire_ni1liiO_dataout;
	wire	wire_ni1lili_dataout;
	wire	wire_ni1lill_dataout;
	wire	wire_ni1lilO_dataout;
	wire	wire_ni1liOi_dataout;
	wire	wire_ni1liOl_dataout;
	wire	wire_ni1liOO_dataout;
	wire	wire_ni1ll0i_dataout;
	wire	wire_ni1ll0l_dataout;
	wire	wire_ni1ll0O_dataout;
	wire	wire_ni1ll1i_dataout;
	wire	wire_ni1ll1l_dataout;
	wire	wire_ni1ll1O_dataout;
	wire	wire_ni1llii_dataout;
	wire	wire_ni1llil_dataout;
	wire	wire_ni1lliO_dataout;
	wire	wire_ni1llli_dataout;
	wire	wire_ni1llll_dataout;
	wire	wire_ni1lllO_dataout;
	wire	wire_ni1llOi_dataout;
	wire	wire_ni1llOl_dataout;
	wire	wire_ni1llOO_dataout;
	wire	wire_ni1lO0i_dataout;
	wire	wire_ni1lO0l_dataout;
	wire	wire_ni1lO0O_dataout;
	wire	wire_ni1lO1i_dataout;
	wire	wire_ni1lO1l_dataout;
	wire	wire_ni1lO1O_dataout;
	wire	wire_ni1lOii_dataout;
	wire	wire_ni1lOil_dataout;
	wire	wire_ni1lOiO_dataout;
	wire	wire_ni1lOli_dataout;
	wire	wire_ni1lOll_dataout;
	wire	wire_ni1lOlO_dataout;
	wire	wire_ni1lOOi_dataout;
	wire	wire_ni1lOOl_dataout;
	wire	wire_ni1lOOO_dataout;
	wire	wire_ni1O00i_dataout;
	wire	wire_ni1O00l_dataout;
	wire	wire_ni1O00O_dataout;
	wire	wire_ni1O01i_dataout;
	wire	wire_ni1O01l_dataout;
	wire	wire_ni1O01O_dataout;
	wire	wire_ni1O0ii_dataout;
	wire	wire_ni1O0il_dataout;
	wire	wire_ni1O0iO_dataout;
	wire	wire_ni1O0li_dataout;
	wire	wire_ni1O0ll_dataout;
	wire	wire_ni1O0lO_dataout;
	wire	wire_ni1O0Oi_dataout;
	wire	wire_ni1O0Ol_dataout;
	wire	wire_ni1O0OO_dataout;
	wire	wire_ni1O10i_dataout;
	wire	wire_ni1O10l_dataout;
	wire	wire_ni1O10O_dataout;
	wire	wire_ni1O11i_dataout;
	wire	wire_ni1O11l_dataout;
	wire	wire_ni1O11O_dataout;
	wire	wire_ni1O1ii_dataout;
	wire	wire_ni1O1il_dataout;
	wire	wire_ni1O1iO_dataout;
	wire	wire_ni1O1li_dataout;
	wire	wire_ni1O1ll_dataout;
	wire	wire_ni1O1lO_dataout;
	wire	wire_ni1O1Oi_dataout;
	wire	wire_ni1O1Ol_dataout;
	wire	wire_ni1O1OO_dataout;
	wire	wire_ni1Oi0i_dataout;
	wire	wire_ni1Oi0l_dataout;
	wire	wire_ni1Oi0O_dataout;
	wire	wire_ni1Oi1i_dataout;
	wire	wire_ni1Oi1l_dataout;
	wire	wire_ni1Oi1O_dataout;
	wire	wire_ni1Oiii_dataout;
	wire	wire_ni1Oiil_dataout;
	wire	wire_ni1OiiO_dataout;
	wire	wire_ni1Oili_dataout;
	wire	wire_ni1Oill_dataout;
	wire	wire_ni1OilO_dataout;
	wire	wire_ni1OiOi_dataout;
	wire	wire_ni1OiOl_dataout;
	wire	wire_ni1OiOO_dataout;
	wire	wire_ni1Ol0i_dataout;
	wire	wire_ni1Ol0l_dataout;
	wire	wire_ni1Ol0O_dataout;
	wire	wire_ni1Ol1i_dataout;
	wire	wire_ni1Ol1l_dataout;
	wire	wire_ni1Ol1O_dataout;
	wire	wire_ni1Olii_dataout;
	wire	wire_ni1Olil_dataout;
	wire	wire_ni1OliO_dataout;
	wire	wire_ni1Olli_dataout;
	wire	wire_ni1Olll_dataout;
	wire	wire_ni1OllO_dataout;
	wire	wire_ni1OlOi_dataout;
	wire	wire_ni1OlOl_dataout;
	wire	wire_ni1OlOO_dataout;
	wire	wire_ni1OO0i_dataout;
	wire	wire_ni1OO0l_dataout;
	wire	wire_ni1OO0O_dataout;
	wire	wire_ni1OO1i_dataout;
	wire	wire_ni1OO1l_dataout;
	wire	wire_ni1OO1O_dataout;
	wire	wire_ni1OOii_dataout;
	wire	wire_ni1OOil_dataout;
	wire	wire_ni1OOiO_dataout;
	wire	wire_ni1OOli_dataout;
	wire	wire_ni1OOll_dataout;
	wire	wire_ni1OOlO_dataout;
	wire	wire_ni1OOOi_dataout;
	wire	wire_ni1OOOl_dataout;
	wire	wire_ni1OOOO_dataout;
	wire	wire_nii001i_dataout;
	wire	wire_nii00ll_dataout;
	wire	wire_nii00lO_dataout;
	wire	wire_nii00Oi_dataout;
	wire	wire_nii00Ol_dataout;
	wire	wire_nii00OO_dataout;
	wire	wire_nii011i_dataout;
	wire	wire_nii01ll_dataout;
	wire	wire_nii01lO_dataout;
	wire	wire_nii01Oi_dataout;
	wire	wire_nii01Ol_dataout;
	wire	wire_nii01OO_dataout;
	wire	wire_nii1OOi_dataout;
	wire	wire_nii1OOl_dataout;
	wire	wire_nii1OOO_dataout;
	wire	wire_niiiO0i_dataout;
	wire	wire_niiiO0l_dataout;
	wire	wire_niiiO0O_dataout;
	wire	wire_niiiO1i_dataout;
	wire	wire_niiiO1l_dataout;
	wire	wire_niiiO1O_dataout;
	wire	wire_niiiOii_dataout;
	wire	wire_niiiOil_dataout;
	wire	wire_niiiOiO_dataout;
	wire	wire_niiiOli_dataout;
	wire	wire_niiiOll_dataout;
	wire	wire_niiiOlO_dataout;
	wire	wire_niiiOOi_dataout;
	wire	wire_niiiOOl_dataout;
	wire	wire_niiiOOO_dataout;
	wire	wire_niil00i_dataout;
	wire	wire_niil00l_dataout;
	wire	wire_niil00O_dataout;
	wire	wire_niil01i_dataout;
	wire	wire_niil01l_dataout;
	wire	wire_niil01O_dataout;
	wire	wire_niil0ii_dataout;
	wire	wire_niil0il_dataout;
	wire	wire_niil0iO_dataout;
	wire	wire_niil0li_dataout;
	wire	wire_niil0ll_dataout;
	wire	wire_niil0lO_dataout;
	wire	wire_niil0Oi_dataout;
	wire	wire_niil0Ol_dataout;
	wire	wire_niil0OO_dataout;
	wire	wire_niil10i_dataout;
	wire	wire_niil10l_dataout;
	wire	wire_niil10O_dataout;
	wire	wire_niil11i_dataout;
	wire	wire_niil11l_dataout;
	wire	wire_niil11O_dataout;
	wire	wire_niil1ii_dataout;
	wire	wire_niil1il_dataout;
	wire	wire_niil1iO_dataout;
	wire	wire_niil1li_dataout;
	wire	wire_niil1ll_dataout;
	wire	wire_niil1lO_dataout;
	wire	wire_niil1Oi_dataout;
	wire	wire_niil1Ol_dataout;
	wire	wire_niil1OO_dataout;
	wire	wire_niili0i_dataout;
	wire	wire_niili0l_dataout;
	wire	wire_niili0O_dataout;
	wire	wire_niili1i_dataout;
	wire	wire_niili1l_dataout;
	wire	wire_niili1O_dataout;
	wire	wire_niiliii_dataout;
	wire	wire_niiliOi_dataout;
	wire	wire_niiliOl_dataout;
	wire	wire_niiliOO_dataout;
	wire	wire_niill0i_dataout;
	wire	wire_niill0l_dataout;
	wire	wire_niill0O_dataout;
	wire	wire_niill1i_dataout;
	wire	wire_niill1l_dataout;
	wire	wire_niill1O_dataout;
	wire	wire_niillii_dataout;
	wire	wire_niillil_dataout;
	wire	wire_niilliO_dataout;
	wire	wire_niillli_dataout;
	wire	wire_niillll_dataout;
	wire	wire_niilllO_dataout;
	wire	wire_niillOi_dataout;
	wire	wire_niillOl_dataout;
	wire	wire_niillOO_dataout;
	wire	wire_niilO0i_dataout;
	wire	wire_niilO0l_dataout;
	wire	wire_niilO0O_dataout;
	wire	wire_niilO1i_dataout;
	wire	wire_niilO1l_dataout;
	wire	wire_niilO1O_dataout;
	wire	wire_niilOii_dataout;
	wire	wire_niilOil_dataout;
	wire	wire_niilOiO_dataout;
	wire	wire_niilOli_dataout;
	wire	wire_niilOll_dataout;
	wire	wire_niilOlO_dataout;
	wire	wire_niilOOi_dataout;
	wire	wire_niilOOl_dataout;
	wire	wire_niilOOO_dataout;
	wire	wire_niiO00i_dataout;
	wire	wire_niiO01i_dataout;
	wire	wire_niiO01l_dataout;
	wire	wire_niiO01O_dataout;
	wire	wire_niiO0iO_dataout;
	wire	wire_niiO0li_dataout;
	wire	wire_niiO0ll_dataout;
	wire	wire_niiO0lO_dataout;
	wire	wire_niiO0Oi_dataout;
	wire	wire_niiO0Ol_dataout;
	wire	wire_niiO0OO_dataout;
	wire	wire_niiO10i_dataout;
	wire	wire_niiO10l_dataout;
	wire	wire_niiO10O_dataout;
	wire	wire_niiO11i_dataout;
	wire	wire_niiO11l_dataout;
	wire	wire_niiO11O_dataout;
	wire	wire_niiO1ii_dataout;
	wire	wire_niiO1il_dataout;
	wire	wire_niiO1iO_dataout;
	wire	wire_niiO1li_dataout;
	wire	wire_niiO1ll_dataout;
	wire	wire_niiO1lO_dataout;
	wire	wire_niiO1Oi_dataout;
	wire	wire_niiO1Ol_dataout;
	wire	wire_niiO1OO_dataout;
	wire	wire_niiOi0i_dataout;
	wire	wire_niiOi0l_dataout;
	wire	wire_niiOi0O_dataout;
	wire	wire_niiOi1i_dataout;
	wire	wire_niiOi1l_dataout;
	wire	wire_niiOi1O_dataout;
	wire	wire_niiOiii_dataout;
	wire	wire_niiOiil_dataout;
	wire	wire_niiOiiO_dataout;
	wire	wire_niiOili_dataout;
	wire	wire_niiOill_dataout;
	wire	wire_niiOilO_dataout;
	wire	wire_niiOiOi_dataout;
	wire	wire_niiOiOl_dataout;
	wire	wire_niiOiOO_dataout;
	wire	wire_niiOl0i_dataout;
	wire	wire_niiOl0l_dataout;
	wire	wire_niiOl0O_dataout;
	wire	wire_niiOl1i_dataout;
	wire	wire_niiOl1l_dataout;
	wire	wire_niiOl1O_dataout;
	wire	wire_niiOlii_dataout;
	wire	wire_niiOlil_dataout;
	wire	wire_niiOliO_dataout;
	wire	wire_niiOlli_dataout;
	wire	wire_niiOlll_dataout;
	wire	wire_niiOllO_dataout;
	wire	wire_niiOlOi_dataout;
	wire	wire_niiOlOl_dataout;
	wire	wire_niiOlOO_dataout;
	wire	wire_niiOO0i_dataout;
	wire	wire_niiOO0l_dataout;
	wire	wire_niiOO0O_dataout;
	wire	wire_niiOO1i_dataout;
	wire	wire_niiOO1l_dataout;
	wire	wire_niiOO1O_dataout;
	wire	wire_niiOOii_dataout;
	wire	wire_niiOOil_dataout;
	wire	wire_niiOOiO_dataout;
	wire	wire_niiOOli_dataout;
	wire	wire_niiOOll_dataout;
	wire	wire_niiOOlO_dataout;
	wire	wire_niiOOOi_dataout;
	wire	wire_niiOOOl_dataout;
	wire	wire_niiOOOO_dataout;
	wire	wire_nil0O0i_dataout;
	wire	wire_nil0O0l_dataout;
	wire	wire_nil0O0O_dataout;
	wire	wire_nil0O1O_dataout;
	wire	wire_nil0Oii_dataout;
	wire	wire_nil0Oil_dataout;
	wire	wire_nil0OiO_dataout;
	wire	wire_nil0Oli_dataout;
	wire	wire_nil0Oll_dataout;
	wire	wire_nil0OlO_dataout;
	wire	wire_nil0OOi_dataout;
	wire	wire_nil0OOl_dataout;
	wire	wire_nil0OOO_dataout;
	wire	wire_nil101i_dataout;
	wire	wire_nil101l_dataout;
	wire	wire_nil10Oi_dataout;
	wire	wire_nil10Ol_dataout;
	wire	wire_nil10OO_dataout;
	wire	wire_nil1i1i_dataout;
	wire	wire_nil1i1l_dataout;
	wire	wire_nili00i_dataout;
	wire	wire_nili00l_dataout;
	wire	wire_nili00O_dataout;
	wire	wire_nili01i_dataout;
	wire	wire_nili01l_dataout;
	wire	wire_nili01O_dataout;
	wire	wire_nili0ii_dataout;
	wire	wire_nili0il_dataout;
	wire	wire_nili0iO_dataout;
	wire	wire_nili0li_dataout;
	wire	wire_nili0ll_dataout;
	wire	wire_nili0lO_dataout;
	wire	wire_nili0Oi_dataout;
	wire	wire_nili0Ol_dataout;
	wire	wire_nili0OO_dataout;
	wire	wire_nili10i_dataout;
	wire	wire_nili10l_dataout;
	wire	wire_nili10O_dataout;
	wire	wire_nili11i_dataout;
	wire	wire_nili11l_dataout;
	wire	wire_nili11O_dataout;
	wire	wire_nili1ii_dataout;
	wire	wire_nili1il_dataout;
	wire	wire_nili1iO_dataout;
	wire	wire_nili1li_dataout;
	wire	wire_nili1ll_dataout;
	wire	wire_nili1lO_dataout;
	wire	wire_nili1Oi_dataout;
	wire	wire_nili1Ol_dataout;
	wire	wire_nili1OO_dataout;
	wire	wire_nilii0i_dataout;
	wire	wire_nilii0l_dataout;
	wire	wire_nilii0O_dataout;
	wire	wire_nilii1i_dataout;
	wire	wire_nilii1l_dataout;
	wire	wire_nilii1O_dataout;
	wire	wire_niliiii_dataout;
	wire	wire_niliiil_dataout;
	wire	wire_niliiiO_dataout;
	wire	wire_niliiOO_dataout;
	wire	wire_nilil0i_dataout;
	wire	wire_nilil0l_dataout;
	wire	wire_nilil0O_dataout;
	wire	wire_nilil1i_dataout;
	wire	wire_nilil1l_dataout;
	wire	wire_nilil1O_dataout;
	wire	wire_nililii_dataout;
	wire	wire_nililil_dataout;
	wire	wire_nililiO_dataout;
	wire	wire_nililli_dataout;
	wire	wire_nililll_dataout;
	wire	wire_nilillO_dataout;
	wire	wire_nililOi_dataout;
	wire	wire_nililOl_dataout;
	wire	wire_nililOO_dataout;
	wire	wire_niliO0i_dataout;
	wire	wire_niliO0l_dataout;
	wire	wire_niliO0O_dataout;
	wire	wire_niliO1i_dataout;
	wire	wire_niliO1l_dataout;
	wire	wire_niliO1O_dataout;
	wire	wire_niliOii_dataout;
	wire	wire_niliOil_dataout;
	wire	wire_niliOiO_dataout;
	wire	wire_niliOli_dataout;
	wire	wire_niliOll_dataout;
	wire	wire_niliOlO_dataout;
	wire	wire_niliOOi_dataout;
	wire	wire_niliOOl_dataout;
	wire	wire_niliOOO_dataout;
	wire	wire_nill00i_dataout;
	wire	wire_nill00l_dataout;
	wire	wire_nill00O_dataout;
	wire	wire_nill01i_dataout;
	wire	wire_nill01l_dataout;
	wire	wire_nill01O_dataout;
	wire	wire_nill0ll_dataout;
	wire	wire_nill0lO_dataout;
	wire	wire_nill0Oi_dataout;
	wire	wire_nill0Ol_dataout;
	wire	wire_nill0OO_dataout;
	wire	wire_nill10i_dataout;
	wire	wire_nill10l_dataout;
	wire	wire_nill10O_dataout;
	wire	wire_nill11i_dataout;
	wire	wire_nill11l_dataout;
	wire	wire_nill11O_dataout;
	wire	wire_nill1ii_dataout;
	wire	wire_nill1il_dataout;
	wire	wire_nill1iO_dataout;
	wire	wire_nill1li_dataout;
	wire	wire_nill1ll_dataout;
	wire	wire_nill1lO_dataout;
	wire	wire_nill1Oi_dataout;
	wire	wire_nill1Ol_dataout;
	wire	wire_nill1OO_dataout;
	wire	wire_nilli0i_dataout;
	wire	wire_nilli0l_dataout;
	wire	wire_nilli0O_dataout;
	wire	wire_nilli1i_dataout;
	wire	wire_nilli1l_dataout;
	wire	wire_nilli1O_dataout;
	wire	wire_nilliii_dataout;
	wire	wire_nilliil_dataout;
	wire	wire_nilliiO_dataout;
	wire	wire_nillili_dataout;
	wire	wire_nillill_dataout;
	wire	wire_nillilO_dataout;
	wire	wire_nilliOi_dataout;
	wire	wire_nilliOl_dataout;
	wire	wire_nilliOO_dataout;
	wire	wire_nilll0i_dataout;
	wire	wire_nilll0l_dataout;
	wire	wire_nilll0O_dataout;
	wire	wire_nilll1i_dataout;
	wire	wire_nilll1l_dataout;
	wire	wire_nilll1O_dataout;
	wire	wire_nilllii_dataout;
	wire	wire_nilllil_dataout;
	wire	wire_nillliO_dataout;
	wire	wire_nilllli_dataout;
	wire	wire_nilllll_dataout;
	wire	wire_nillllO_dataout;
	wire	wire_nilllOi_dataout;
	wire	wire_nilllOl_dataout;
	wire	wire_nilllOO_dataout;
	wire	wire_nillO0i_dataout;
	wire	wire_nillO0l_dataout;
	wire	wire_nillO0O_dataout;
	wire	wire_nillO1i_dataout;
	wire	wire_nillO1l_dataout;
	wire	wire_nillO1O_dataout;
	wire	wire_nillOii_dataout;
	wire	wire_nillOil_dataout;
	wire	wire_nillOiO_dataout;
	wire	wire_nillOli_dataout;
	wire	wire_nillOll_dataout;
	wire	wire_nillOlO_dataout;
	wire	wire_nillOOi_dataout;
	wire	wire_nillOOl_dataout;
	wire	wire_nillOOO_dataout;
	wire	wire_nilO00i_dataout;
	wire	wire_nilO00O_dataout;
	wire	wire_nilO01O_dataout;
	wire	wire_nilO0ii_dataout;
	wire	wire_nilO0il_dataout;
	wire	wire_nilO0lO_dataout;
	wire	wire_nilO0OO_dataout;
	wire	wire_nilO11i_dataout;
	wire	wire_nilO11l_dataout;
	wire	wire_nilOi1l_dataout;
	wire	wire_nilOiOO_dataout;
	wire	wire_nilOl0i_dataout;
	wire	wire_nilOl1i_dataout;
	wire	wire_nilOl1l_dataout;
	wire	wire_nilOl1O_dataout;
	wire	wire_niO00li_dataout;
	wire	wire_niO00ll_dataout;
	wire	wire_niO010i_dataout;
	wire	wire_niO010l_dataout;
	wire	wire_niO010O_dataout;
	wire	wire_niO011i_dataout;
	wire	wire_niO011l_dataout;
	wire	wire_niO011O_dataout;
	wire	wire_niO01ii_dataout;
	wire	wire_niO01il_dataout;
	wire	wire_niO01iO_dataout;
	wire	wire_niO100i_dataout;
	wire	wire_niO100l_dataout;
	wire	wire_niO100O_dataout;
	wire	wire_niO101i_dataout;
	wire	wire_niO101l_dataout;
	wire	wire_niO101O_dataout;
	wire	wire_niO10ii_dataout;
	wire	wire_niO10il_dataout;
	wire	wire_niO10iO_dataout;
	wire	wire_niO10li_dataout;
	wire	wire_niO10ll_dataout;
	wire	wire_niO10lO_dataout;
	wire	wire_niO10Oi_dataout;
	wire	wire_niO10Ol_dataout;
	wire	wire_niO10OO_dataout;
	wire	wire_niO1i0i_dataout;
	wire	wire_niO1i0l_dataout;
	wire	wire_niO1i1i_dataout;
	wire	wire_niO1i1l_dataout;
	wire	wire_niO1i1O_dataout;
	wire	wire_niO1ill_dataout;
	wire	wire_niO1ilO_dataout;
	wire	wire_niO1iOi_dataout;
	wire	wire_niO1iOl_dataout;
	wire	wire_niO1iOO_dataout;
	wire	wire_niO1l0i_dataout;
	wire	wire_niO1l0l_dataout;
	wire	wire_niO1l0O_dataout;
	wire	wire_niO1l1i_dataout;
	wire	wire_niO1l1l_dataout;
	wire	wire_niO1l1O_dataout;
	wire	wire_niO1lii_dataout;
	wire	wire_niO1lil_dataout;
	wire	wire_niO1liO_dataout;
	wire	wire_niO1lli_dataout;
	wire	wire_niO1lll_dataout;
	wire	wire_niO1llO_dataout;
	wire	wire_niO1lOi_dataout;
	wire	wire_niO1lOl_dataout;
	wire	wire_niO1lOO_dataout;
	wire	wire_niO1O0l_dataout;
	wire	wire_niO1O0O_dataout;
	wire	wire_niO1Oii_dataout;
	wire	wire_niO1Oil_dataout;
	wire	wire_niO1OiO_dataout;
	wire	wire_niO1Oli_dataout;
	wire	wire_niO1Oll_dataout;
	wire	wire_niO1OlO_dataout;
	wire	wire_niO1OOi_dataout;
	wire	wire_niO1OOl_dataout;
	wire	wire_niO1OOO_dataout;
	wire	wire_niOiOil_dataout;
	wire	wire_niOiOiO_dataout;
	wire	wire_niOl00i_dataout;
	wire	wire_niOl00l_dataout;
	wire	wire_niOl00O_dataout;
	wire	wire_niOl01i_dataout;
	wire	wire_niOl01l_dataout;
	wire	wire_niOl01O_dataout;
	wire	wire_niOl0ii_dataout;
	wire	wire_niOl10l_dataout;
	wire	wire_niOl10O_dataout;
	wire	wire_niOl1ii_dataout;
	wire	wire_niOl1il_dataout;
	wire	wire_niOl1iO_dataout;
	wire	wire_niOl1li_dataout;
	wire	wire_niOl1ll_dataout;
	wire	wire_niOl1lO_dataout;
	wire	wire_niOl1Oi_dataout;
	wire	wire_niOl1Ol_dataout;
	wire	wire_niOl1OO_dataout;
	wire	wire_nl0i00i_dataout;
	wire	wire_nl0i00l_dataout;
	wire	wire_nl0i00O_dataout;
	wire	wire_nl0i01i_dataout;
	wire	wire_nl0i01l_dataout;
	wire	wire_nl0i01O_dataout;
	wire	wire_nl0i0ii_dataout;
	wire	wire_nl0i1OO_dataout;
	wire	wire_nl0iill_dataout;
	wire	wire_nl0iilO_dataout;
	wire	wire_nl0iiOi_dataout;
	wire	wire_nl0iiOl_dataout;
	wire	wire_nl0iiOO_dataout;
	wire	wire_nl0il0i_dataout;
	wire	wire_nl0il0l_dataout;
	wire	wire_nl0il1i_dataout;
	wire	wire_nl0il1l_dataout;
	wire	wire_nl0il1O_dataout;
	wire	wire_nl0iO0i_dataout;
	wire	wire_nl0iO0l_dataout;
	wire	wire_nl0iO0O_dataout;
	wire	wire_nl0iOii_dataout;
	wire	wire_nl0iOil_dataout;
	wire	wire_nl0iOiO_dataout;
	wire	wire_nl0iOli_dataout;
	wire	wire_nl0iOll_dataout;
	wire	wire_nl0iOlO_dataout;
	wire	wire_nl0iOOi_dataout;
	wire	wire_nl0l01i_dataout;
	wire	wire_nl0l01l_dataout;
	wire	wire_nl0O10i_dataout;
	wire	wire_nl0O10l_dataout;
	wire	wire_nl0O10O_dataout;
	wire	wire_nl0O11i_dataout;
	wire	wire_nl0O11l_dataout;
	wire	wire_nl0O11O_dataout;
	wire	wire_nl0O1ii_dataout;
	wire	wire_nl0O1il_dataout;
	wire	wire_nl0O1iO_dataout;
	wire	wire_nl0O1li_dataout;
	wire	wire_nl0O1ll_dataout;
	wire	wire_nl1lO0l_dataout;
	wire	wire_nl1lO0O_dataout;
	wire	wire_nl1lOii_dataout;
	wire	wire_nl1lOil_dataout;
	wire	wire_nl1lOiO_dataout;
	wire	wire_nl1lOli_dataout;
	wire	wire_nl1lOll_dataout;
	wire	wire_nl1lOlO_dataout;
	wire	wire_nl1O0ii_dataout;
	wire	wire_nl1O0il_dataout;
	wire	wire_nl1O0iO_dataout;
	wire	wire_nl1O0li_dataout;
	wire	wire_nl1O0ll_dataout;
	wire	wire_nl1O0lO_dataout;
	wire	wire_nl1O0Oi_dataout;
	wire	wire_nl1O0Ol_dataout;
	wire	wire_nl1O0OO_dataout;
	wire  [1:0]   wire_ni010Ol_o;
	wire  [2:0]   wire_ni01i1l_o;
	wire  [1:0]   wire_ni01iOO_o;
	wire  [2:0]   wire_ni01l0i_o;
	wire  [1:0]   wire_ni01lOO_o;
	wire  [2:0]   wire_ni01O1O_o;
	wire  [0:0]   wire_ni0Oiil_o;
	wire  [1:0]   wire_ni0Oili_o;
	wire  [6:0]   wire_nii001l_o;
	wire  [4:0]   wire_nii011l_o;
	wire  [10:0]   wire_niOO1lO_o;
	wire  [8:0]   wire_niOOi0l_o;
	wire  [8:0]   wire_nl0i0il_o;
	wire  [10:0]   wire_nl0il0O_o;
	wire  [10:0]   wire_nl0iOOl_o;
	wire  [3:0]   wire_nl0l01O_o;
	wire  [9:0]   wire_nl0O00O_o;
	wire  [11:0]   wire_nl0O0ii_o;
	wire  [12:0]   wire_nl0O1lO_o;
	wire  [11:0]   wire_nl0O1Oi_o;
	wire  [8:0]   wire_nl0Olil_o;
	wire  [11:0]   wire_nl0OOii_o;
	wire  [18:0]   wire_nl1iOll_o;
	wire  [18:0]   wire_nl1l01O_o;
	wire  [18:0]   wire_nl1l1ii_o;
	wire  [8:0]   wire_nl1lOOi_o;
	wire  [10:0]   wire_nl1Oi1i_o;
	wire  [11:0]   wire_nli110l_o;
	wire  [9:0]   wire_nli110O_o;
	wire  [9:0]   wire_nli11ii_o;
	wire  wire_nii111l_o;
	wire  wire_n011i_o;
	wire  wire_n011l_o;
	wire  wire_n1ilO_o;
	wire  wire_n1iOi_o;
	wire  wire_n1iOl_o;
	wire  wire_n1iOO_o;
	wire  wire_n1l0i_o;
	wire  wire_n1l0l_o;
	wire  wire_n1l0O_o;
	wire  wire_n1l1i_o;
	wire  wire_n1l1l_o;
	wire  wire_n1l1O_o;
	wire  wire_n1lii_o;
	wire  wire_n1lil_o;
	wire  wire_n1liO_o;
	wire  wire_n1lli_o;
	wire  wire_n1lll_o;
	wire  wire_n1llO_o;
	wire  wire_n1lOi_o;
	wire  wire_n1lOl_o;
	wire  wire_n1lOO_o;
	wire  wire_n1O0i_o;
	wire  wire_n1O0l_o;
	wire  wire_n1O0O_o;
	wire  wire_n1O1i_o;
	wire  wire_n1O1l_o;
	wire  wire_n1O1O_o;
	wire  wire_n1Oii_o;
	wire  wire_n1Oil_o;
	wire  wire_n1OiO_o;
	wire  wire_n1Oli_o;
	wire  wire_n1Oll_o;
	wire  wire_n1OlO_o;
	wire  wire_n1OOi_o;
	wire  wire_n1OOl_o;
	wire  wire_n1OOO_o;
	wire  wire_ni00i_o;
	wire  wire_ni00l_o;
	wire  wire_ni00O_o;
	wire  wire_ni01i_o;
	wire  wire_ni01l_o;
	wire  wire_ni01O_o;
	wire  wire_ni0ii_o;
	wire  wire_ni0il_o;
	wire  wire_ni0iO_o;
	wire  wire_ni0li_o;
	wire  wire_ni0ll_o;
	wire  wire_ni0lO_o;
	wire  wire_ni0Oi_o;
	wire  wire_ni0Ol_o;
	wire  wire_ni0OO_o;
	wire  wire_ni10O_o;
	wire  wire_ni1ii_o;
	wire  wire_ni1il_o;
	wire  wire_ni1iO_o;
	wire  wire_ni1li_o;
	wire  wire_ni1ll_o;
	wire  wire_ni1lO_o;
	wire  wire_ni1Oi_o;
	wire  wire_ni1Ol_o;
	wire  wire_ni1OO_o;
	wire  wire_nii0i_o;
	wire  wire_nii0l_o;
	wire  wire_nii0O_o;
	wire  wire_nii1i_o;
	wire  wire_nii1l_o;
	wire  wire_nii1O_o;
	wire  wire_niiii_o;
	wire  wire_niiil_o;
	wire  wire_niiiO_o;
	wire  wire_niili_o;
	wire  wire_niill_o;
	wire  wire_niilO_o;
	wire  wire_niiOi_o;
	wire  wire_niiOl_o;
	wire  wire_niiOO_o;
	wire  wire_nil0i_o;
	wire  wire_nil0l_o;
	wire  wire_nil0O_o;
	wire  wire_nil1i_o;
	wire  wire_nil1l_o;
	wire  wire_nil1O_o;
	wire  wire_nilii_o;
	wire  wire_nilil_o;
	wire  wire_niliO_o;
	wire  wire_nilli_o;
	wire  wire_nilll_o;
	wire  wire_nillO_o;
	wire  wire_nilOi_o;
	wire  wire_nilOl_o;
	wire  wire_nilOO_o;
	wire  wire_niO0i_o;
	wire  wire_niO0l_o;
	wire  wire_niO0O_o;
	wire  wire_niO1i_o;
	wire  wire_niO1l_o;
	wire  wire_niO1O_o;
	wire  wire_niOii_o;
	wire  wire_niOil_o;
	wire  wire_niOiO_o;
	wire  wire_niOli_o;
	wire  wire_niOll_o;
	wire  wire_niOlO_o;
	wire  wire_niOOi_o;
	wire  wire_niOOl_o;
	wire  wire_nlO10O_o;
	wire  wire_nlO1ii_o;
	wire  wire_nlO1il_o;
	wire  wire_nlO1iO_o;
	wire  wire_nlO1li_o;
	wire  wire_nlO1ll_o;
	wire  wire_ni011ii_o;
	wire  wire_ni011Ol_o;
	wire  wire_nii00ii_o;
	wire  wire_nii11iO_o;
	wire  wire_nii1O0O_o;
	wire  wire_nil10iO_o;
	wire  wire_nilOill_o;
	wire  wire_niO0i1l_o;
	wire  wire_niO0ili_o;
	wire  wire_niO0O0O_o;
	wire  wire_niO0Oii_o;
	wire  wire_niO0Oil_o;
	wire  wire_niO0OiO_o;
	wire  wire_niO0Oli_o;
	wire  wire_niO0Oll_o;
	wire  wire_niO0OlO_o;
	wire  wire_niO0OOi_o;
	wire  wire_niO0OOl_o;
	wire  wire_niO0OOO_o;
	wire  wire_niOi00O_o;
	wire  wire_niOi0Oi_o;
	wire  wire_niOi10i_o;
	wire  wire_niOi10l_o;
	wire  wire_niOi10O_o;
	wire  wire_niOi11i_o;
	wire  wire_niOi11l_o;
	wire  wire_niOi11O_o;
	wire  wire_niOi1ii_o;
	wire  wire_niOi1il_o;
	wire  wire_niOi1iO_o;
	wire  wire_niOi1li_o;
	wire  wire_niOi1ll_o;
	wire  wire_niOi1lO_o;
	wire  wire_niOi1Oi_o;
	wire  wire_niOi1Ol_o;
	wire  wire_niOll0O_o;
	wire  wire_niOllii_o;
	wire  wire_niOllil_o;
	wire  wire_niOlliO_o;
	wire  wire_niOllli_o;
	wire  wire_niOllll_o;
	wire  wire_niOlllO_o;
	wire  wire_niOllOi_o;
	wire  wire_niOllOl_o;
	wire  wire_niOllOO_o;
	wire  wire_niOlOOl_o;
	wire  wire_niOO0iO_o;
	wire  wire_niOOlOO_o;
	wire  wire_niOOO0i_o;
	wire  wire_niOOO0l_o;
	wire  wire_niOOO0O_o;
	wire  wire_niOOO1i_o;
	wire  wire_niOOO1l_o;
	wire  wire_niOOO1O_o;
	wire  wire_niOOOii_o;
	wire  wire_niOOOil_o;
	wire  wire_niOOOiO_o;
	wire  wire_niOOOli_o;
	wire  wire_niOOOll_o;
	wire  wire_niOOOlO_o;
	wire  wire_niOOOOi_o;
	wire  wire_niOOOOl_o;
	wire  wire_niOOOOO_o;
	wire  wire_nl000iO_o;
	wire  wire_nl000li_o;
	wire  wire_nl000ll_o;
	wire  wire_nl000lO_o;
	wire  wire_nl000Oi_o;
	wire  wire_nl000Ol_o;
	wire  wire_nl000OO_o;
	wire  wire_nl0010O_o;
	wire  wire_nl00i1i_o;
	wire  wire_nl00i1l_o;
	wire  wire_nl00i1O_o;
	wire  wire_nl010ll_o;
	wire  wire_nl010lO_o;
	wire  wire_nl010Oi_o;
	wire  wire_nl010Ol_o;
	wire  wire_nl0111l_o;
	wire  wire_nl0111O_o;
	wire  wire_nl011lO_o;
	wire  wire_nl011Oi_o;
	wire  wire_nl011Ol_o;
	wire  wire_nl011OO_o;
	wire  wire_nl01lii_o;
	wire  wire_nl01O1i_o;
	wire  wire_nl01Oli_o;
	wire  wire_nl0l00l_o;
	wire  wire_nl0l0li_o;
	wire  wire_nl0llii_o;
	wire  wire_nl0llil_o;
	wire  wire_nl0lliO_o;
	wire  wire_nl0llli_o;
	wire  wire_nl0llll_o;
	wire  wire_nl0lllO_o;
	wire  wire_nl0llOi_o;
	wire  wire_nl0llOl_o;
	wire  wire_nl0llOO_o;
	wire  wire_nl0lO1i_o;
	wire  wire_nl0lO1l_o;
	wire  wire_nl1000O_o;
	wire  wire_nl1010i_o;
	wire  wire_nl1010l_o;
	wire  wire_nl1010O_o;
	wire  wire_nl1011i_o;
	wire  wire_nl1011l_o;
	wire  wire_nl1011O_o;
	wire  wire_nl101ii_o;
	wire  wire_nl101il_o;
	wire  wire_nl101iO_o;
	wire  wire_nl101li_o;
	wire  wire_nl101ll_o;
	wire  wire_nl101lO_o;
	wire  wire_nl101Oi_o;
	wire  wire_nl101Ol_o;
	wire  wire_nl101OO_o;
	wire  wire_nl1110i_o;
	wire  wire_nl1110l_o;
	wire  wire_nl1110O_o;
	wire  wire_nl1111i_o;
	wire  wire_nl1111l_o;
	wire  wire_nl1111O_o;
	wire  wire_nl111ii_o;
	wire  wire_nl111il_o;
	wire  wire_nl111Ol_o;
	wire  wire_nl11Oii_o;
	wire  wire_nl11Oil_o;
	wire  wire_nl11OiO_o;
	wire  wire_nl11Oli_o;
	wire  wire_nl11Oll_o;
	wire  wire_nl11OlO_o;
	wire  wire_nl11OOi_o;
	wire  wire_nl11OOl_o;
	wire  wire_nl11OOO_o;
	wire  wire_nl1l0lO_o;
	wire  wire_nl1l0Oi_o;
	wire  wire_nl1l0Ol_o;
	wire  wire_nl1l0OO_o;
	wire  wire_nl1li0i_o;
	wire  wire_nl1li1i_o;
	wire  wire_nl1li1l_o;
	wire  wire_nl1li1O_o;
	wire  wire_nl1liOi_o;
	wire  wire_nl1liOl_o;
	wire  wire_nl1liOO_o;
	wire  wire_nl1ll0i_o;
	wire  wire_nl1ll0l_o;
	wire  wire_nl1ll1i_o;
	wire  wire_nl1ll1l_o;
	wire  wire_nl1ll1O_o;
	wire  wire_nl1llii_o;
	wire  wire_nl1lliO_o;
	wire  n0OOili;
	wire  n0OOill;
	wire  n0OOilO;
	wire  n0OOiOi;
	wire  n0OOiOl;
	wire  n0OOiOO;
	wire  n0OOl0i;
	wire  n0OOl0l;
	wire  n0OOl0O;
	wire  n0OOl1i;
	wire  n0OOl1l;
	wire  n0OOl1O;
	wire  n0OOlii;
	wire  n0OOlil;
	wire  n0OOliO;
	wire  n0OOlli;
	wire  n0OOlll;
	wire  n0OOllO;
	wire  n0OOlOi;
	wire  n0OOlOl;
	wire  n0OOlOO;
	wire  n0OOO0i;
	wire  n0OOO0l;
	wire  n0OOO0O;
	wire  n0OOO1i;
	wire  n0OOO1l;
	wire  n0OOO1O;
	wire  n0OOOii;
	wire  n0OOOil;
	wire  n0OOOiO;
	wire  n0OOOli;
	wire  n0OOOll;
	wire  n0OOOlO;
	wire  n0OOOOi;
	wire  n0OOOOl;
	wire  n0OOOOO;
	wire  ni1000i;
	wire  ni1000l;
	wire  ni1000O;
	wire  ni1001i;
	wire  ni1001l;
	wire  ni1001O;
	wire  ni100ii;
	wire  ni100il;
	wire  ni100iO;
	wire  ni100li;
	wire  ni100ll;
	wire  ni100lO;
	wire  ni100Oi;
	wire  ni100Ol;
	wire  ni100OO;
	wire  ni1010i;
	wire  ni1010l;
	wire  ni1010O;
	wire  ni1011i;
	wire  ni1011l;
	wire  ni1011O;
	wire  ni101ii;
	wire  ni101il;
	wire  ni101iO;
	wire  ni101li;
	wire  ni101ll;
	wire  ni101lO;
	wire  ni101Oi;
	wire  ni101Ol;
	wire  ni101OO;
	wire  ni10i0i;
	wire  ni10i0l;
	wire  ni10i0O;
	wire  ni10i1i;
	wire  ni10i1l;
	wire  ni10i1O;
	wire  ni10iii;
	wire  ni10iil;
	wire  ni10iiO;
	wire  ni10ili;
	wire  ni10ill;
	wire  ni10ilO;
	wire  ni10iOi;
	wire  ni10iOl;
	wire  ni10iOO;
	wire  ni10l0i;
	wire  ni10l0l;
	wire  ni10l0O;
	wire  ni10l1i;
	wire  ni10l1l;
	wire  ni10l1O;
	wire  ni10lii;
	wire  ni10lil;
	wire  ni10liO;
	wire  ni10lli;
	wire  ni10lll;
	wire  ni10llO;
	wire  ni10lOi;
	wire  ni10lOl;
	wire  ni10lOO;
	wire  ni10O0i;
	wire  ni10O0l;
	wire  ni10O0O;
	wire  ni10O1i;
	wire  ni10O1l;
	wire  ni10O1O;
	wire  ni10Oii;
	wire  ni10Oil;
	wire  ni10OiO;
	wire  ni10Oli;
	wire  ni10Oll;
	wire  ni10OlO;
	wire  ni10OOi;
	wire  ni10OOl;
	wire  ni10OOO;
	wire  ni1100i;
	wire  ni1100l;
	wire  ni1100O;
	wire  ni1101i;
	wire  ni1101l;
	wire  ni1101O;
	wire  ni110ii;
	wire  ni110il;
	wire  ni110iO;
	wire  ni110li;
	wire  ni110ll;
	wire  ni110lO;
	wire  ni110Oi;
	wire  ni110Ol;
	wire  ni110OO;
	wire  ni1110i;
	wire  ni1110l;
	wire  ni1110O;
	wire  ni1111i;
	wire  ni1111l;
	wire  ni1111O;
	wire  ni111ii;
	wire  ni111il;
	wire  ni111iO;
	wire  ni111li;
	wire  ni111ll;
	wire  ni111lO;
	wire  ni111Oi;
	wire  ni111Ol;
	wire  ni111OO;
	wire  ni11i0i;
	wire  ni11i0l;
	wire  ni11i0O;
	wire  ni11i1i;
	wire  ni11i1l;
	wire  ni11i1O;
	wire  ni11iii;
	wire  ni11iil;
	wire  ni11iiO;
	wire  ni11ili;
	wire  ni11ill;
	wire  ni11ilO;
	wire  ni11iOi;
	wire  ni11iOl;
	wire  ni11iOO;
	wire  ni11l0i;
	wire  ni11l0l;
	wire  ni11l0O;
	wire  ni11l1i;
	wire  ni11l1l;
	wire  ni11l1O;
	wire  ni11lii;
	wire  ni11lil;
	wire  ni11liO;
	wire  ni11lli;
	wire  ni11lll;
	wire  ni11llO;
	wire  ni11lOi;
	wire  ni11lOl;
	wire  ni11lOO;
	wire  ni11O0i;
	wire  ni11O0l;
	wire  ni11O0O;
	wire  ni11O1i;
	wire  ni11O1l;
	wire  ni11O1O;
	wire  ni11Oii;
	wire  ni11Oil;
	wire  ni11OiO;
	wire  ni11Oli;
	wire  ni11Oll;
	wire  ni11OlO;
	wire  ni11OOi;
	wire  ni11OOl;
	wire  ni11OOO;
	wire  ni1i00i;
	wire  ni1i01l;
	wire  ni1i0ii;
	wire  ni1i0li;
	wire  ni1i0lO;
	wire  ni1i0OO;
	wire  ni1i10i;
	wire  ni1i10l;
	wire  ni1i11i;
	wire  ni1i11l;
	wire  ni1i11O;
	wire  ni1i1il;
	wire  ni1i1iO;
	wire  ni1i1lO;
	wire  ni1i1OO;
	wire  ni1ii0i;
	wire  ni1ii0l;
	wire  ni1ii0O;
	wire  ni1ii1l;
	wire  ni1iiii;
	wire  ni1iiil;
	wire  ni1iiiO;
	wire  ni1iili;
	wire  ni1iilO;
	wire  ni1iiOi;
	wire  ni1iiOl;
	wire  ni1iiOO;
	wire  ni1il1i;
	wire  ni1il1l;
	wire  ni1iOli;

	altmult_add   nl1Oi1O
	( 
	.chainout_sat_overflow(),
	.clock0(clock),
	.dataa({nl1O1li, nl1O1il, nl1O1ii, nl1O10O, nl1O10l, nl1O10i, nl1O11O, nl1O11l, nl1O11i}),
	.datab({1'b0, nli0l0l, nli0l1O, nli0l1l, nli0l1i, nli0iOO, nli0iOl, nli0iOi, nli0ilO}),
	.ena0(((~ ni1iili) & ((n010l | nl1Oiil) | nl1Oi0i))),
	.mult0_is_saturated(),
	.mult1_is_saturated(),
	.mult2_is_saturated(),
	.mult3_is_saturated(),
	.overflow(),
	.result(wire_nl1Oi1O_result),
	.scanouta(),
	.scanoutb(),
	.signa(1'b0),
	.signb(1'b0),
	.accum_sload(),
	.aclr0(),
	.aclr1(),
	.aclr2(),
	.aclr3(),
	.addnsub1(),
	.addnsub1_round(),
	.addnsub3(),
	.addnsub3_round(),
	.chainin(),
	.chainout_round(),
	.chainout_saturate(),
	.clock1(),
	.clock2(),
	.clock3(),
	.coefsel0(),
	.coefsel1(),
	.coefsel2(),
	.coefsel3(),
	.datac(),
	.ena1(),
	.ena2(),
	.ena3(),
	.mult01_round(),
	.mult01_saturation(),
	.mult23_round(),
	.mult23_saturation(),
	.output_round(),
	.output_saturate(),
	.rotate(),
	.scanina(),
	.scaninb(),
	.shift_right(),
	.sourcea(),
	.sourceb(),
	.zero_chainout(),
	.zero_loopback()
	);
	defparam
		nl1Oi1O.accum_direction = "ADD",
		nl1Oi1O.accum_sload_aclr = "ACLR3",
		nl1Oi1O.accum_sload_pipeline_aclr = "ACLR3",
		nl1Oi1O.accum_sload_pipeline_register = "CLOCK0",
		nl1Oi1O.accum_sload_register = "CLOCK0",
		nl1Oi1O.accumulator = "NO",
		nl1Oi1O.adder1_rounding = "NO",
		nl1Oi1O.adder3_rounding = "NO",
		nl1Oi1O.addnsub1_round_aclr = "ACLR3",
		nl1Oi1O.addnsub1_round_pipeline_aclr = "ACLR3",
		nl1Oi1O.addnsub1_round_pipeline_register = "CLOCK0",
		nl1Oi1O.addnsub1_round_register = "CLOCK0",
		nl1Oi1O.addnsub3_round_aclr = "ACLR3",
		nl1Oi1O.addnsub3_round_pipeline_aclr = "ACLR3",
		nl1Oi1O.addnsub3_round_pipeline_register = "CLOCK0",
		nl1Oi1O.addnsub3_round_register = "CLOCK0",
		nl1Oi1O.addnsub_multiplier_aclr1 = "ACLR3",
		nl1Oi1O.addnsub_multiplier_aclr3 = "ACLR3",
		nl1Oi1O.addnsub_multiplier_pipeline_aclr1 = "ACLR3",
		nl1Oi1O.addnsub_multiplier_pipeline_aclr3 = "ACLR3",
		nl1Oi1O.addnsub_multiplier_pipeline_register1 = "UNREGISTERED",
		nl1Oi1O.addnsub_multiplier_pipeline_register3 = "UNREGISTERED",
		nl1Oi1O.addnsub_multiplier_register1 = "CLOCK0",
		nl1Oi1O.addnsub_multiplier_register3 = "CLOCK0",
		nl1Oi1O.chainout_aclr = "ACLR3",
		nl1Oi1O.chainout_adder = "NO",
		nl1Oi1O.chainout_register = "CLOCK0",
		nl1Oi1O.chainout_round_aclr = "ACLR3",
		nl1Oi1O.chainout_round_output_aclr = "ACLR3",
		nl1Oi1O.chainout_round_output_register = "CLOCK0",
		nl1Oi1O.chainout_round_pipeline_aclr = "ACLR3",
		nl1Oi1O.chainout_round_pipeline_register = "CLOCK0",
		nl1Oi1O.chainout_round_register = "CLOCK0",
		nl1Oi1O.chainout_rounding = "NO",
		nl1Oi1O.chainout_saturate_aclr = "ACLR3",
		nl1Oi1O.chainout_saturate_output_aclr = "ACLR3",
		nl1Oi1O.chainout_saturate_output_register = "CLOCK0",
		nl1Oi1O.chainout_saturate_pipeline_aclr = "ACLR3",
		nl1Oi1O.chainout_saturate_pipeline_register = "CLOCK0",
		nl1Oi1O.chainout_saturate_register = "CLOCK0",
		nl1Oi1O.chainout_saturation = "NO",
		nl1Oi1O.coef0_0 = 0,
		nl1Oi1O.coef0_1 = 0,
		nl1Oi1O.coef0_2 = 0,
		nl1Oi1O.coef0_3 = 0,
		nl1Oi1O.coef0_4 = 0,
		nl1Oi1O.coef0_5 = 0,
		nl1Oi1O.coef0_6 = 0,
		nl1Oi1O.coef0_7 = 0,
		nl1Oi1O.coef1_0 = 0,
		nl1Oi1O.coef1_1 = 0,
		nl1Oi1O.coef1_2 = 0,
		nl1Oi1O.coef1_3 = 0,
		nl1Oi1O.coef1_4 = 0,
		nl1Oi1O.coef1_5 = 0,
		nl1Oi1O.coef1_6 = 0,
		nl1Oi1O.coef1_7 = 0,
		nl1Oi1O.coef2_0 = 0,
		nl1Oi1O.coef2_1 = 0,
		nl1Oi1O.coef2_2 = 0,
		nl1Oi1O.coef2_3 = 0,
		nl1Oi1O.coef2_4 = 0,
		nl1Oi1O.coef2_5 = 0,
		nl1Oi1O.coef2_6 = 0,
		nl1Oi1O.coef2_7 = 0,
		nl1Oi1O.coef3_0 = 0,
		nl1Oi1O.coef3_1 = 0,
		nl1Oi1O.coef3_2 = 0,
		nl1Oi1O.coef3_3 = 0,
		nl1Oi1O.coef3_4 = 0,
		nl1Oi1O.coef3_5 = 0,
		nl1Oi1O.coef3_6 = 0,
		nl1Oi1O.coef3_7 = 0,
		nl1Oi1O.coefsel0_aclr = "ACLR0",
		nl1Oi1O.coefsel0_register = "CLOCK0",
		nl1Oi1O.coefsel1_aclr = "ACLR0",
		nl1Oi1O.coefsel1_register = "CLOCK0",
		nl1Oi1O.coefsel2_aclr = "ACLR0",
		nl1Oi1O.coefsel2_register = "CLOCK0",
		nl1Oi1O.coefsel3_aclr = "ACLR0",
		nl1Oi1O.coefsel3_register = "CLOCK0",
		nl1Oi1O.dsp_block_balancing = "AUTO",
		nl1Oi1O.extra_latency = 0,
		nl1Oi1O.input_aclr_a0 = "ACLR3",
		nl1Oi1O.input_aclr_a1 = "ACLR3",
		nl1Oi1O.input_aclr_a2 = "ACLR3",
		nl1Oi1O.input_aclr_a3 = "ACLR3",
		nl1Oi1O.input_aclr_b0 = "ACLR3",
		nl1Oi1O.input_aclr_b1 = "ACLR3",
		nl1Oi1O.input_aclr_b2 = "ACLR3",
		nl1Oi1O.input_aclr_b3 = "ACLR3",
		nl1Oi1O.input_aclr_c0 = "ACLR0",
		nl1Oi1O.input_register_a0 = "CLOCK0",
		nl1Oi1O.input_register_a1 = "CLOCK0",
		nl1Oi1O.input_register_a2 = "CLOCK0",
		nl1Oi1O.input_register_a3 = "CLOCK0",
		nl1Oi1O.input_register_b0 = "CLOCK0",
		nl1Oi1O.input_register_b1 = "CLOCK0",
		nl1Oi1O.input_register_b2 = "CLOCK0",
		nl1Oi1O.input_register_b3 = "CLOCK0",
		nl1Oi1O.input_register_c0 = "CLOCK0",
		nl1Oi1O.input_source_a0 = "DATAA",
		nl1Oi1O.input_source_a1 = "DATAA",
		nl1Oi1O.input_source_a2 = "DATAA",
		nl1Oi1O.input_source_a3 = "DATAA",
		nl1Oi1O.input_source_b0 = "DATAB",
		nl1Oi1O.input_source_b1 = "DATAB",
		nl1Oi1O.input_source_b2 = "DATAB",
		nl1Oi1O.input_source_b3 = "DATAB",
		nl1Oi1O.intended_device_family = "Cyclone III",
		nl1Oi1O.loadconst_value = 64,
		nl1Oi1O.mult01_round_aclr = "ACLR3",
		nl1Oi1O.mult01_round_register = "CLOCK0",
		nl1Oi1O.mult01_saturation_aclr = "ACLR2",
		nl1Oi1O.mult01_saturation_register = "CLOCK0",
		nl1Oi1O.mult23_round_aclr = "ACLR3",
		nl1Oi1O.mult23_round_register = "CLOCK0",
		nl1Oi1O.mult23_saturation_aclr = "ACLR3",
		nl1Oi1O.mult23_saturation_register = "CLOCK0",
		nl1Oi1O.multiplier01_rounding = "NO",
		nl1Oi1O.multiplier01_saturation = "NO",
		nl1Oi1O.multiplier1_direction = "ADD",
		nl1Oi1O.multiplier23_rounding = "NO",
		nl1Oi1O.multiplier23_saturation = "NO",
		nl1Oi1O.multiplier3_direction = "ADD",
		nl1Oi1O.multiplier_aclr0 = "ACLR3",
		nl1Oi1O.multiplier_aclr1 = "ACLR3",
		nl1Oi1O.multiplier_aclr2 = "ACLR3",
		nl1Oi1O.multiplier_aclr3 = "ACLR3",
		nl1Oi1O.multiplier_register0 = "CLOCK0",
		nl1Oi1O.multiplier_register1 = "CLOCK0",
		nl1Oi1O.multiplier_register2 = "CLOCK0",
		nl1Oi1O.multiplier_register3 = "CLOCK0",
		nl1Oi1O.number_of_multipliers = 1,
		nl1Oi1O.output_aclr = "ACLR0",
		nl1Oi1O.output_register = "CLOCK0",
		nl1Oi1O.output_round_aclr = "ACLR3",
		nl1Oi1O.output_round_pipeline_aclr = "ACLR3",
		nl1Oi1O.output_round_pipeline_register = "CLOCK0",
		nl1Oi1O.output_round_register = "CLOCK0",
		nl1Oi1O.output_round_type = "NEAREST_INTEGER",
		nl1Oi1O.output_rounding = "NO",
		nl1Oi1O.output_saturate_aclr = "ACLR3",
		nl1Oi1O.output_saturate_pipeline_aclr = "ACLR3",
		nl1Oi1O.output_saturate_pipeline_register = "CLOCK0",
		nl1Oi1O.output_saturate_register = "CLOCK0",
		nl1Oi1O.output_saturate_type = "ASYMMETRIC",
		nl1Oi1O.output_saturation = "NO",
		nl1Oi1O.port_addnsub1 = "PORT_UNUSED",
		nl1Oi1O.port_addnsub3 = "PORT_UNUSED",
		nl1Oi1O.port_chainout_sat_is_overflow = "PORT_UNUSED",
		nl1Oi1O.port_output_is_overflow = "PORT_UNUSED",
		nl1Oi1O.port_signa = "PORT_CONNECTIVITY",
		nl1Oi1O.port_signb = "PORT_CONNECTIVITY",
		nl1Oi1O.preadder_direction_0 = "ADD",
		nl1Oi1O.preadder_direction_1 = "ADD",
		nl1Oi1O.preadder_direction_2 = "ADD",
		nl1Oi1O.preadder_direction_3 = "ADD",
		nl1Oi1O.preadder_mode = "SIMPLE",
		nl1Oi1O.representation_a = "UNSIGNED",
		nl1Oi1O.representation_b = "UNSIGNED",
		nl1Oi1O.rotate_aclr = "ACLR3",
		nl1Oi1O.rotate_output_aclr = "ACLR3",
		nl1Oi1O.rotate_output_register = "CLOCK0",
		nl1Oi1O.rotate_pipeline_aclr = "ACLR3",
		nl1Oi1O.rotate_pipeline_register = "CLOCK0",
		nl1Oi1O.rotate_register = "CLOCK0",
		nl1Oi1O.scanouta_aclr = "ACLR3",
		nl1Oi1O.scanouta_register = "UNREGISTERED",
		nl1Oi1O.shift_mode = "NO",
		nl1Oi1O.shift_right_aclr = "ACLR3",
		nl1Oi1O.shift_right_output_aclr = "ACLR3",
		nl1Oi1O.shift_right_output_register = "CLOCK0",
		nl1Oi1O.shift_right_pipeline_aclr = "ACLR3",
		nl1Oi1O.shift_right_pipeline_register = "CLOCK0",
		nl1Oi1O.shift_right_register = "CLOCK0",
		nl1Oi1O.signed_aclr_a = "ACLR3",
		nl1Oi1O.signed_aclr_b = "ACLR3",
		nl1Oi1O.signed_pipeline_aclr_a = "ACLR3",
		nl1Oi1O.signed_pipeline_aclr_b = "ACLR3",
		nl1Oi1O.signed_pipeline_register_a = "UNREGISTERED",
		nl1Oi1O.signed_pipeline_register_b = "UNREGISTERED",
		nl1Oi1O.signed_register_a = "CLOCK0",
		nl1Oi1O.signed_register_b = "CLOCK0",
		nl1Oi1O.systolic_aclr1 = "ACLR0",
		nl1Oi1O.systolic_aclr3 = "ACLR0",
		nl1Oi1O.systolic_delay1 = "UNREGISTERED",
		nl1Oi1O.systolic_delay3 = "UNREGISTERED",
		nl1Oi1O.width_a = 9,
		nl1Oi1O.width_b = 9,
		nl1Oi1O.width_c = 22,
		nl1Oi1O.width_chainin = 1,
		nl1Oi1O.width_coef = 18,
		nl1Oi1O.width_msb = 17,
		nl1Oi1O.width_result = 18,
		nl1Oi1O.width_saturate_sign = 1,
		nl1Oi1O.zero_chainout_output_aclr = "ACLR3",
		nl1Oi1O.zero_chainout_output_register = "CLOCK0",
		nl1Oi1O.zero_loopback_aclr = "ACLR3",
		nl1Oi1O.zero_loopback_output_aclr = "ACLR3",
		nl1Oi1O.zero_loopback_output_register = "CLOCK0",
		nl1Oi1O.zero_loopback_pipeline_aclr = "ACLR3",
		nl1Oi1O.zero_loopback_pipeline_register = "CLOCK0",
		nl1Oi1O.zero_loopback_register = "CLOCK0";
	altmult_add   nl1OiiO
	( 
	.chainout_sat_overflow(),
	.clock0(clock),
	.dataa({nl1O1li, nl1O1il, nl1O1ii, nl1O10O, nl1O10l, nl1O10i, nl1O11O, nl1O11l, nl1O11i}),
	.datab({1'b0, nli0lOO, nli0lOi, nli0llO, nli0lll, nli0lli, nli0liO, nli0lil, nli0lii}),
	.ena0(((~ ni1iili) & ((n010l | nl1OiOl) | nl1Oili))),
	.mult0_is_saturated(),
	.mult1_is_saturated(),
	.mult2_is_saturated(),
	.mult3_is_saturated(),
	.overflow(),
	.result(wire_nl1OiiO_result),
	.scanouta(),
	.scanoutb(),
	.signa(1'b0),
	.signb(1'b0),
	.accum_sload(),
	.aclr0(),
	.aclr1(),
	.aclr2(),
	.aclr3(),
	.addnsub1(),
	.addnsub1_round(),
	.addnsub3(),
	.addnsub3_round(),
	.chainin(),
	.chainout_round(),
	.chainout_saturate(),
	.clock1(),
	.clock2(),
	.clock3(),
	.coefsel0(),
	.coefsel1(),
	.coefsel2(),
	.coefsel3(),
	.datac(),
	.ena1(),
	.ena2(),
	.ena3(),
	.mult01_round(),
	.mult01_saturation(),
	.mult23_round(),
	.mult23_saturation(),
	.output_round(),
	.output_saturate(),
	.rotate(),
	.scanina(),
	.scaninb(),
	.shift_right(),
	.sourcea(),
	.sourceb(),
	.zero_chainout(),
	.zero_loopback()
	);
	defparam
		nl1OiiO.accum_direction = "ADD",
		nl1OiiO.accum_sload_aclr = "ACLR3",
		nl1OiiO.accum_sload_pipeline_aclr = "ACLR3",
		nl1OiiO.accum_sload_pipeline_register = "CLOCK0",
		nl1OiiO.accum_sload_register = "CLOCK0",
		nl1OiiO.accumulator = "NO",
		nl1OiiO.adder1_rounding = "NO",
		nl1OiiO.adder3_rounding = "NO",
		nl1OiiO.addnsub1_round_aclr = "ACLR3",
		nl1OiiO.addnsub1_round_pipeline_aclr = "ACLR3",
		nl1OiiO.addnsub1_round_pipeline_register = "CLOCK0",
		nl1OiiO.addnsub1_round_register = "CLOCK0",
		nl1OiiO.addnsub3_round_aclr = "ACLR3",
		nl1OiiO.addnsub3_round_pipeline_aclr = "ACLR3",
		nl1OiiO.addnsub3_round_pipeline_register = "CLOCK0",
		nl1OiiO.addnsub3_round_register = "CLOCK0",
		nl1OiiO.addnsub_multiplier_aclr1 = "ACLR3",
		nl1OiiO.addnsub_multiplier_aclr3 = "ACLR3",
		nl1OiiO.addnsub_multiplier_pipeline_aclr1 = "ACLR3",
		nl1OiiO.addnsub_multiplier_pipeline_aclr3 = "ACLR3",
		nl1OiiO.addnsub_multiplier_pipeline_register1 = "UNREGISTERED",
		nl1OiiO.addnsub_multiplier_pipeline_register3 = "UNREGISTERED",
		nl1OiiO.addnsub_multiplier_register1 = "CLOCK0",
		nl1OiiO.addnsub_multiplier_register3 = "CLOCK0",
		nl1OiiO.chainout_aclr = "ACLR3",
		nl1OiiO.chainout_adder = "NO",
		nl1OiiO.chainout_register = "CLOCK0",
		nl1OiiO.chainout_round_aclr = "ACLR3",
		nl1OiiO.chainout_round_output_aclr = "ACLR3",
		nl1OiiO.chainout_round_output_register = "CLOCK0",
		nl1OiiO.chainout_round_pipeline_aclr = "ACLR3",
		nl1OiiO.chainout_round_pipeline_register = "CLOCK0",
		nl1OiiO.chainout_round_register = "CLOCK0",
		nl1OiiO.chainout_rounding = "NO",
		nl1OiiO.chainout_saturate_aclr = "ACLR3",
		nl1OiiO.chainout_saturate_output_aclr = "ACLR3",
		nl1OiiO.chainout_saturate_output_register = "CLOCK0",
		nl1OiiO.chainout_saturate_pipeline_aclr = "ACLR3",
		nl1OiiO.chainout_saturate_pipeline_register = "CLOCK0",
		nl1OiiO.chainout_saturate_register = "CLOCK0",
		nl1OiiO.chainout_saturation = "NO",
		nl1OiiO.coef0_0 = 0,
		nl1OiiO.coef0_1 = 0,
		nl1OiiO.coef0_2 = 0,
		nl1OiiO.coef0_3 = 0,
		nl1OiiO.coef0_4 = 0,
		nl1OiiO.coef0_5 = 0,
		nl1OiiO.coef0_6 = 0,
		nl1OiiO.coef0_7 = 0,
		nl1OiiO.coef1_0 = 0,
		nl1OiiO.coef1_1 = 0,
		nl1OiiO.coef1_2 = 0,
		nl1OiiO.coef1_3 = 0,
		nl1OiiO.coef1_4 = 0,
		nl1OiiO.coef1_5 = 0,
		nl1OiiO.coef1_6 = 0,
		nl1OiiO.coef1_7 = 0,
		nl1OiiO.coef2_0 = 0,
		nl1OiiO.coef2_1 = 0,
		nl1OiiO.coef2_2 = 0,
		nl1OiiO.coef2_3 = 0,
		nl1OiiO.coef2_4 = 0,
		nl1OiiO.coef2_5 = 0,
		nl1OiiO.coef2_6 = 0,
		nl1OiiO.coef2_7 = 0,
		nl1OiiO.coef3_0 = 0,
		nl1OiiO.coef3_1 = 0,
		nl1OiiO.coef3_2 = 0,
		nl1OiiO.coef3_3 = 0,
		nl1OiiO.coef3_4 = 0,
		nl1OiiO.coef3_5 = 0,
		nl1OiiO.coef3_6 = 0,
		nl1OiiO.coef3_7 = 0,
		nl1OiiO.coefsel0_aclr = "ACLR0",
		nl1OiiO.coefsel0_register = "CLOCK0",
		nl1OiiO.coefsel1_aclr = "ACLR0",
		nl1OiiO.coefsel1_register = "CLOCK0",
		nl1OiiO.coefsel2_aclr = "ACLR0",
		nl1OiiO.coefsel2_register = "CLOCK0",
		nl1OiiO.coefsel3_aclr = "ACLR0",
		nl1OiiO.coefsel3_register = "CLOCK0",
		nl1OiiO.dsp_block_balancing = "AUTO",
		nl1OiiO.extra_latency = 0,
		nl1OiiO.input_aclr_a0 = "ACLR3",
		nl1OiiO.input_aclr_a1 = "ACLR3",
		nl1OiiO.input_aclr_a2 = "ACLR3",
		nl1OiiO.input_aclr_a3 = "ACLR3",
		nl1OiiO.input_aclr_b0 = "ACLR3",
		nl1OiiO.input_aclr_b1 = "ACLR3",
		nl1OiiO.input_aclr_b2 = "ACLR3",
		nl1OiiO.input_aclr_b3 = "ACLR3",
		nl1OiiO.input_aclr_c0 = "ACLR0",
		nl1OiiO.input_register_a0 = "CLOCK0",
		nl1OiiO.input_register_a1 = "CLOCK0",
		nl1OiiO.input_register_a2 = "CLOCK0",
		nl1OiiO.input_register_a3 = "CLOCK0",
		nl1OiiO.input_register_b0 = "CLOCK0",
		nl1OiiO.input_register_b1 = "CLOCK0",
		nl1OiiO.input_register_b2 = "CLOCK0",
		nl1OiiO.input_register_b3 = "CLOCK0",
		nl1OiiO.input_register_c0 = "CLOCK0",
		nl1OiiO.input_source_a0 = "DATAA",
		nl1OiiO.input_source_a1 = "DATAA",
		nl1OiiO.input_source_a2 = "DATAA",
		nl1OiiO.input_source_a3 = "DATAA",
		nl1OiiO.input_source_b0 = "DATAB",
		nl1OiiO.input_source_b1 = "DATAB",
		nl1OiiO.input_source_b2 = "DATAB",
		nl1OiiO.input_source_b3 = "DATAB",
		nl1OiiO.intended_device_family = "Cyclone III",
		nl1OiiO.loadconst_value = 64,
		nl1OiiO.mult01_round_aclr = "ACLR3",
		nl1OiiO.mult01_round_register = "CLOCK0",
		nl1OiiO.mult01_saturation_aclr = "ACLR2",
		nl1OiiO.mult01_saturation_register = "CLOCK0",
		nl1OiiO.mult23_round_aclr = "ACLR3",
		nl1OiiO.mult23_round_register = "CLOCK0",
		nl1OiiO.mult23_saturation_aclr = "ACLR3",
		nl1OiiO.mult23_saturation_register = "CLOCK0",
		nl1OiiO.multiplier01_rounding = "NO",
		nl1OiiO.multiplier01_saturation = "NO",
		nl1OiiO.multiplier1_direction = "ADD",
		nl1OiiO.multiplier23_rounding = "NO",
		nl1OiiO.multiplier23_saturation = "NO",
		nl1OiiO.multiplier3_direction = "ADD",
		nl1OiiO.multiplier_aclr0 = "ACLR3",
		nl1OiiO.multiplier_aclr1 = "ACLR3",
		nl1OiiO.multiplier_aclr2 = "ACLR3",
		nl1OiiO.multiplier_aclr3 = "ACLR3",
		nl1OiiO.multiplier_register0 = "CLOCK0",
		nl1OiiO.multiplier_register1 = "CLOCK0",
		nl1OiiO.multiplier_register2 = "CLOCK0",
		nl1OiiO.multiplier_register3 = "CLOCK0",
		nl1OiiO.number_of_multipliers = 1,
		nl1OiiO.output_aclr = "ACLR0",
		nl1OiiO.output_register = "CLOCK0",
		nl1OiiO.output_round_aclr = "ACLR3",
		nl1OiiO.output_round_pipeline_aclr = "ACLR3",
		nl1OiiO.output_round_pipeline_register = "CLOCK0",
		nl1OiiO.output_round_register = "CLOCK0",
		nl1OiiO.output_round_type = "NEAREST_INTEGER",
		nl1OiiO.output_rounding = "NO",
		nl1OiiO.output_saturate_aclr = "ACLR3",
		nl1OiiO.output_saturate_pipeline_aclr = "ACLR3",
		nl1OiiO.output_saturate_pipeline_register = "CLOCK0",
		nl1OiiO.output_saturate_register = "CLOCK0",
		nl1OiiO.output_saturate_type = "ASYMMETRIC",
		nl1OiiO.output_saturation = "NO",
		nl1OiiO.port_addnsub1 = "PORT_UNUSED",
		nl1OiiO.port_addnsub3 = "PORT_UNUSED",
		nl1OiiO.port_chainout_sat_is_overflow = "PORT_UNUSED",
		nl1OiiO.port_output_is_overflow = "PORT_UNUSED",
		nl1OiiO.port_signa = "PORT_CONNECTIVITY",
		nl1OiiO.port_signb = "PORT_CONNECTIVITY",
		nl1OiiO.preadder_direction_0 = "ADD",
		nl1OiiO.preadder_direction_1 = "ADD",
		nl1OiiO.preadder_direction_2 = "ADD",
		nl1OiiO.preadder_direction_3 = "ADD",
		nl1OiiO.preadder_mode = "SIMPLE",
		nl1OiiO.representation_a = "UNSIGNED",
		nl1OiiO.representation_b = "UNSIGNED",
		nl1OiiO.rotate_aclr = "ACLR3",
		nl1OiiO.rotate_output_aclr = "ACLR3",
		nl1OiiO.rotate_output_register = "CLOCK0",
		nl1OiiO.rotate_pipeline_aclr = "ACLR3",
		nl1OiiO.rotate_pipeline_register = "CLOCK0",
		nl1OiiO.rotate_register = "CLOCK0",
		nl1OiiO.scanouta_aclr = "ACLR3",
		nl1OiiO.scanouta_register = "UNREGISTERED",
		nl1OiiO.shift_mode = "NO",
		nl1OiiO.shift_right_aclr = "ACLR3",
		nl1OiiO.shift_right_output_aclr = "ACLR3",
		nl1OiiO.shift_right_output_register = "CLOCK0",
		nl1OiiO.shift_right_pipeline_aclr = "ACLR3",
		nl1OiiO.shift_right_pipeline_register = "CLOCK0",
		nl1OiiO.shift_right_register = "CLOCK0",
		nl1OiiO.signed_aclr_a = "ACLR3",
		nl1OiiO.signed_aclr_b = "ACLR3",
		nl1OiiO.signed_pipeline_aclr_a = "ACLR3",
		nl1OiiO.signed_pipeline_aclr_b = "ACLR3",
		nl1OiiO.signed_pipeline_register_a = "UNREGISTERED",
		nl1OiiO.signed_pipeline_register_b = "UNREGISTERED",
		nl1OiiO.signed_register_a = "CLOCK0",
		nl1OiiO.signed_register_b = "CLOCK0",
		nl1OiiO.systolic_aclr1 = "ACLR0",
		nl1OiiO.systolic_aclr3 = "ACLR0",
		nl1OiiO.systolic_delay1 = "UNREGISTERED",
		nl1OiiO.systolic_delay3 = "UNREGISTERED",
		nl1OiiO.width_a = 9,
		nl1OiiO.width_b = 9,
		nl1OiiO.width_c = 22,
		nl1OiiO.width_chainin = 1,
		nl1OiiO.width_coef = 18,
		nl1OiiO.width_msb = 17,
		nl1OiiO.width_result = 18,
		nl1OiiO.width_saturate_sign = 1,
		nl1OiiO.zero_chainout_output_aclr = "ACLR3",
		nl1OiiO.zero_chainout_output_register = "CLOCK0",
		nl1OiiO.zero_loopback_aclr = "ACLR3",
		nl1OiiO.zero_loopback_output_aclr = "ACLR3",
		nl1OiiO.zero_loopback_output_register = "CLOCK0",
		nl1OiiO.zero_loopback_pipeline_aclr = "ACLR3",
		nl1OiiO.zero_loopback_pipeline_register = "CLOCK0",
		nl1OiiO.zero_loopback_register = "CLOCK0";
	altmult_add   nl1OiOO
	( 
	.chainout_sat_overflow(),
	.clock0(clock),
	.dataa({nl1O1li, nl1O1il, nl1O1ii, nl1O10O, nl1O10l, nl1O10i, nl1O11O, nl1O11l, nl1O11i}),
	.datab({1'b0, nli0ili, nli0iil, nli0iii, nli0i0O, nli0i0l, nli0i0i, nli0i1O, nli0i1l}),
	.ena0(((~ ni1iili) & ((n010l | nl1Ol0l) | nl1Ol1i))),
	.mult0_is_saturated(),
	.mult1_is_saturated(),
	.mult2_is_saturated(),
	.mult3_is_saturated(),
	.overflow(),
	.result(wire_nl1OiOO_result),
	.scanouta(),
	.scanoutb(),
	.signa(1'b0),
	.signb(1'b0),
	.accum_sload(),
	.aclr0(),
	.aclr1(),
	.aclr2(),
	.aclr3(),
	.addnsub1(),
	.addnsub1_round(),
	.addnsub3(),
	.addnsub3_round(),
	.chainin(),
	.chainout_round(),
	.chainout_saturate(),
	.clock1(),
	.clock2(),
	.clock3(),
	.coefsel0(),
	.coefsel1(),
	.coefsel2(),
	.coefsel3(),
	.datac(),
	.ena1(),
	.ena2(),
	.ena3(),
	.mult01_round(),
	.mult01_saturation(),
	.mult23_round(),
	.mult23_saturation(),
	.output_round(),
	.output_saturate(),
	.rotate(),
	.scanina(),
	.scaninb(),
	.shift_right(),
	.sourcea(),
	.sourceb(),
	.zero_chainout(),
	.zero_loopback()
	);
	defparam
		nl1OiOO.accum_direction = "ADD",
		nl1OiOO.accum_sload_aclr = "ACLR3",
		nl1OiOO.accum_sload_pipeline_aclr = "ACLR3",
		nl1OiOO.accum_sload_pipeline_register = "CLOCK0",
		nl1OiOO.accum_sload_register = "CLOCK0",
		nl1OiOO.accumulator = "NO",
		nl1OiOO.adder1_rounding = "NO",
		nl1OiOO.adder3_rounding = "NO",
		nl1OiOO.addnsub1_round_aclr = "ACLR3",
		nl1OiOO.addnsub1_round_pipeline_aclr = "ACLR3",
		nl1OiOO.addnsub1_round_pipeline_register = "CLOCK0",
		nl1OiOO.addnsub1_round_register = "CLOCK0",
		nl1OiOO.addnsub3_round_aclr = "ACLR3",
		nl1OiOO.addnsub3_round_pipeline_aclr = "ACLR3",
		nl1OiOO.addnsub3_round_pipeline_register = "CLOCK0",
		nl1OiOO.addnsub3_round_register = "CLOCK0",
		nl1OiOO.addnsub_multiplier_aclr1 = "ACLR3",
		nl1OiOO.addnsub_multiplier_aclr3 = "ACLR3",
		nl1OiOO.addnsub_multiplier_pipeline_aclr1 = "ACLR3",
		nl1OiOO.addnsub_multiplier_pipeline_aclr3 = "ACLR3",
		nl1OiOO.addnsub_multiplier_pipeline_register1 = "UNREGISTERED",
		nl1OiOO.addnsub_multiplier_pipeline_register3 = "UNREGISTERED",
		nl1OiOO.addnsub_multiplier_register1 = "CLOCK0",
		nl1OiOO.addnsub_multiplier_register3 = "CLOCK0",
		nl1OiOO.chainout_aclr = "ACLR3",
		nl1OiOO.chainout_adder = "NO",
		nl1OiOO.chainout_register = "CLOCK0",
		nl1OiOO.chainout_round_aclr = "ACLR3",
		nl1OiOO.chainout_round_output_aclr = "ACLR3",
		nl1OiOO.chainout_round_output_register = "CLOCK0",
		nl1OiOO.chainout_round_pipeline_aclr = "ACLR3",
		nl1OiOO.chainout_round_pipeline_register = "CLOCK0",
		nl1OiOO.chainout_round_register = "CLOCK0",
		nl1OiOO.chainout_rounding = "NO",
		nl1OiOO.chainout_saturate_aclr = "ACLR3",
		nl1OiOO.chainout_saturate_output_aclr = "ACLR3",
		nl1OiOO.chainout_saturate_output_register = "CLOCK0",
		nl1OiOO.chainout_saturate_pipeline_aclr = "ACLR3",
		nl1OiOO.chainout_saturate_pipeline_register = "CLOCK0",
		nl1OiOO.chainout_saturate_register = "CLOCK0",
		nl1OiOO.chainout_saturation = "NO",
		nl1OiOO.coef0_0 = 0,
		nl1OiOO.coef0_1 = 0,
		nl1OiOO.coef0_2 = 0,
		nl1OiOO.coef0_3 = 0,
		nl1OiOO.coef0_4 = 0,
		nl1OiOO.coef0_5 = 0,
		nl1OiOO.coef0_6 = 0,
		nl1OiOO.coef0_7 = 0,
		nl1OiOO.coef1_0 = 0,
		nl1OiOO.coef1_1 = 0,
		nl1OiOO.coef1_2 = 0,
		nl1OiOO.coef1_3 = 0,
		nl1OiOO.coef1_4 = 0,
		nl1OiOO.coef1_5 = 0,
		nl1OiOO.coef1_6 = 0,
		nl1OiOO.coef1_7 = 0,
		nl1OiOO.coef2_0 = 0,
		nl1OiOO.coef2_1 = 0,
		nl1OiOO.coef2_2 = 0,
		nl1OiOO.coef2_3 = 0,
		nl1OiOO.coef2_4 = 0,
		nl1OiOO.coef2_5 = 0,
		nl1OiOO.coef2_6 = 0,
		nl1OiOO.coef2_7 = 0,
		nl1OiOO.coef3_0 = 0,
		nl1OiOO.coef3_1 = 0,
		nl1OiOO.coef3_2 = 0,
		nl1OiOO.coef3_3 = 0,
		nl1OiOO.coef3_4 = 0,
		nl1OiOO.coef3_5 = 0,
		nl1OiOO.coef3_6 = 0,
		nl1OiOO.coef3_7 = 0,
		nl1OiOO.coefsel0_aclr = "ACLR0",
		nl1OiOO.coefsel0_register = "CLOCK0",
		nl1OiOO.coefsel1_aclr = "ACLR0",
		nl1OiOO.coefsel1_register = "CLOCK0",
		nl1OiOO.coefsel2_aclr = "ACLR0",
		nl1OiOO.coefsel2_register = "CLOCK0",
		nl1OiOO.coefsel3_aclr = "ACLR0",
		nl1OiOO.coefsel3_register = "CLOCK0",
		nl1OiOO.dsp_block_balancing = "AUTO",
		nl1OiOO.extra_latency = 0,
		nl1OiOO.input_aclr_a0 = "ACLR3",
		nl1OiOO.input_aclr_a1 = "ACLR3",
		nl1OiOO.input_aclr_a2 = "ACLR3",
		nl1OiOO.input_aclr_a3 = "ACLR3",
		nl1OiOO.input_aclr_b0 = "ACLR3",
		nl1OiOO.input_aclr_b1 = "ACLR3",
		nl1OiOO.input_aclr_b2 = "ACLR3",
		nl1OiOO.input_aclr_b3 = "ACLR3",
		nl1OiOO.input_aclr_c0 = "ACLR0",
		nl1OiOO.input_register_a0 = "CLOCK0",
		nl1OiOO.input_register_a1 = "CLOCK0",
		nl1OiOO.input_register_a2 = "CLOCK0",
		nl1OiOO.input_register_a3 = "CLOCK0",
		nl1OiOO.input_register_b0 = "CLOCK0",
		nl1OiOO.input_register_b1 = "CLOCK0",
		nl1OiOO.input_register_b2 = "CLOCK0",
		nl1OiOO.input_register_b3 = "CLOCK0",
		nl1OiOO.input_register_c0 = "CLOCK0",
		nl1OiOO.input_source_a0 = "DATAA",
		nl1OiOO.input_source_a1 = "DATAA",
		nl1OiOO.input_source_a2 = "DATAA",
		nl1OiOO.input_source_a3 = "DATAA",
		nl1OiOO.input_source_b0 = "DATAB",
		nl1OiOO.input_source_b1 = "DATAB",
		nl1OiOO.input_source_b2 = "DATAB",
		nl1OiOO.input_source_b3 = "DATAB",
		nl1OiOO.intended_device_family = "Cyclone III",
		nl1OiOO.loadconst_value = 64,
		nl1OiOO.mult01_round_aclr = "ACLR3",
		nl1OiOO.mult01_round_register = "CLOCK0",
		nl1OiOO.mult01_saturation_aclr = "ACLR2",
		nl1OiOO.mult01_saturation_register = "CLOCK0",
		nl1OiOO.mult23_round_aclr = "ACLR3",
		nl1OiOO.mult23_round_register = "CLOCK0",
		nl1OiOO.mult23_saturation_aclr = "ACLR3",
		nl1OiOO.mult23_saturation_register = "CLOCK0",
		nl1OiOO.multiplier01_rounding = "NO",
		nl1OiOO.multiplier01_saturation = "NO",
		nl1OiOO.multiplier1_direction = "ADD",
		nl1OiOO.multiplier23_rounding = "NO",
		nl1OiOO.multiplier23_saturation = "NO",
		nl1OiOO.multiplier3_direction = "ADD",
		nl1OiOO.multiplier_aclr0 = "ACLR3",
		nl1OiOO.multiplier_aclr1 = "ACLR3",
		nl1OiOO.multiplier_aclr2 = "ACLR3",
		nl1OiOO.multiplier_aclr3 = "ACLR3",
		nl1OiOO.multiplier_register0 = "CLOCK0",
		nl1OiOO.multiplier_register1 = "CLOCK0",
		nl1OiOO.multiplier_register2 = "CLOCK0",
		nl1OiOO.multiplier_register3 = "CLOCK0",
		nl1OiOO.number_of_multipliers = 1,
		nl1OiOO.output_aclr = "ACLR0",
		nl1OiOO.output_register = "CLOCK0",
		nl1OiOO.output_round_aclr = "ACLR3",
		nl1OiOO.output_round_pipeline_aclr = "ACLR3",
		nl1OiOO.output_round_pipeline_register = "CLOCK0",
		nl1OiOO.output_round_register = "CLOCK0",
		nl1OiOO.output_round_type = "NEAREST_INTEGER",
		nl1OiOO.output_rounding = "NO",
		nl1OiOO.output_saturate_aclr = "ACLR3",
		nl1OiOO.output_saturate_pipeline_aclr = "ACLR3",
		nl1OiOO.output_saturate_pipeline_register = "CLOCK0",
		nl1OiOO.output_saturate_register = "CLOCK0",
		nl1OiOO.output_saturate_type = "ASYMMETRIC",
		nl1OiOO.output_saturation = "NO",
		nl1OiOO.port_addnsub1 = "PORT_UNUSED",
		nl1OiOO.port_addnsub3 = "PORT_UNUSED",
		nl1OiOO.port_chainout_sat_is_overflow = "PORT_UNUSED",
		nl1OiOO.port_output_is_overflow = "PORT_UNUSED",
		nl1OiOO.port_signa = "PORT_CONNECTIVITY",
		nl1OiOO.port_signb = "PORT_CONNECTIVITY",
		nl1OiOO.preadder_direction_0 = "ADD",
		nl1OiOO.preadder_direction_1 = "ADD",
		nl1OiOO.preadder_direction_2 = "ADD",
		nl1OiOO.preadder_direction_3 = "ADD",
		nl1OiOO.preadder_mode = "SIMPLE",
		nl1OiOO.representation_a = "UNSIGNED",
		nl1OiOO.representation_b = "UNSIGNED",
		nl1OiOO.rotate_aclr = "ACLR3",
		nl1OiOO.rotate_output_aclr = "ACLR3",
		nl1OiOO.rotate_output_register = "CLOCK0",
		nl1OiOO.rotate_pipeline_aclr = "ACLR3",
		nl1OiOO.rotate_pipeline_register = "CLOCK0",
		nl1OiOO.rotate_register = "CLOCK0",
		nl1OiOO.scanouta_aclr = "ACLR3",
		nl1OiOO.scanouta_register = "UNREGISTERED",
		nl1OiOO.shift_mode = "NO",
		nl1OiOO.shift_right_aclr = "ACLR3",
		nl1OiOO.shift_right_output_aclr = "ACLR3",
		nl1OiOO.shift_right_output_register = "CLOCK0",
		nl1OiOO.shift_right_pipeline_aclr = "ACLR3",
		nl1OiOO.shift_right_pipeline_register = "CLOCK0",
		nl1OiOO.shift_right_register = "CLOCK0",
		nl1OiOO.signed_aclr_a = "ACLR3",
		nl1OiOO.signed_aclr_b = "ACLR3",
		nl1OiOO.signed_pipeline_aclr_a = "ACLR3",
		nl1OiOO.signed_pipeline_aclr_b = "ACLR3",
		nl1OiOO.signed_pipeline_register_a = "UNREGISTERED",
		nl1OiOO.signed_pipeline_register_b = "UNREGISTERED",
		nl1OiOO.signed_register_a = "CLOCK0",
		nl1OiOO.signed_register_b = "CLOCK0",
		nl1OiOO.systolic_aclr1 = "ACLR0",
		nl1OiOO.systolic_aclr3 = "ACLR0",
		nl1OiOO.systolic_delay1 = "UNREGISTERED",
		nl1OiOO.systolic_delay3 = "UNREGISTERED",
		nl1OiOO.width_a = 9,
		nl1OiOO.width_b = 9,
		nl1OiOO.width_c = 22,
		nl1OiOO.width_chainin = 1,
		nl1OiOO.width_coef = 18,
		nl1OiOO.width_msb = 17,
		nl1OiOO.width_result = 18,
		nl1OiOO.width_saturate_sign = 1,
		nl1OiOO.zero_chainout_output_aclr = "ACLR3",
		nl1OiOO.zero_chainout_output_register = "CLOCK0",
		nl1OiOO.zero_loopback_aclr = "ACLR3",
		nl1OiOO.zero_loopback_output_aclr = "ACLR3",
		nl1OiOO.zero_loopback_output_register = "CLOCK0",
		nl1OiOO.zero_loopback_pipeline_aclr = "ACLR3",
		nl1OiOO.zero_loopback_pipeline_register = "CLOCK0",
		nl1OiOO.zero_loopback_register = "CLOCK0";
	altmult_add   nl1Ol0O
	( 
	.chainout_sat_overflow(),
	.clock0(clock),
	.dataa({nl1O00i, nl1O01O, nl1O01l, nl1O01i, nl1O1OO, nl1O1Ol, nl1O1Oi, nl1O1lO, nl1O00O}),
	.datab({1'b0, nli00OO, nli00Oi, nli00lO, nli00ll, nli00li, nli00iO, nli00il, nli00ii}),
	.ena0(((~ ni1iili) & ((n010l | nl1Olll) | nl1Olii))),
	.mult0_is_saturated(),
	.mult1_is_saturated(),
	.mult2_is_saturated(),
	.mult3_is_saturated(),
	.overflow(),
	.result(wire_nl1Ol0O_result),
	.scanouta(),
	.scanoutb(),
	.signa(1'b0),
	.signb(1'b0),
	.accum_sload(),
	.aclr0(),
	.aclr1(),
	.aclr2(),
	.aclr3(),
	.addnsub1(),
	.addnsub1_round(),
	.addnsub3(),
	.addnsub3_round(),
	.chainin(),
	.chainout_round(),
	.chainout_saturate(),
	.clock1(),
	.clock2(),
	.clock3(),
	.coefsel0(),
	.coefsel1(),
	.coefsel2(),
	.coefsel3(),
	.datac(),
	.ena1(),
	.ena2(),
	.ena3(),
	.mult01_round(),
	.mult01_saturation(),
	.mult23_round(),
	.mult23_saturation(),
	.output_round(),
	.output_saturate(),
	.rotate(),
	.scanina(),
	.scaninb(),
	.shift_right(),
	.sourcea(),
	.sourceb(),
	.zero_chainout(),
	.zero_loopback()
	);
	defparam
		nl1Ol0O.accum_direction = "ADD",
		nl1Ol0O.accum_sload_aclr = "ACLR3",
		nl1Ol0O.accum_sload_pipeline_aclr = "ACLR3",
		nl1Ol0O.accum_sload_pipeline_register = "CLOCK0",
		nl1Ol0O.accum_sload_register = "CLOCK0",
		nl1Ol0O.accumulator = "NO",
		nl1Ol0O.adder1_rounding = "NO",
		nl1Ol0O.adder3_rounding = "NO",
		nl1Ol0O.addnsub1_round_aclr = "ACLR3",
		nl1Ol0O.addnsub1_round_pipeline_aclr = "ACLR3",
		nl1Ol0O.addnsub1_round_pipeline_register = "CLOCK0",
		nl1Ol0O.addnsub1_round_register = "CLOCK0",
		nl1Ol0O.addnsub3_round_aclr = "ACLR3",
		nl1Ol0O.addnsub3_round_pipeline_aclr = "ACLR3",
		nl1Ol0O.addnsub3_round_pipeline_register = "CLOCK0",
		nl1Ol0O.addnsub3_round_register = "CLOCK0",
		nl1Ol0O.addnsub_multiplier_aclr1 = "ACLR3",
		nl1Ol0O.addnsub_multiplier_aclr3 = "ACLR3",
		nl1Ol0O.addnsub_multiplier_pipeline_aclr1 = "ACLR3",
		nl1Ol0O.addnsub_multiplier_pipeline_aclr3 = "ACLR3",
		nl1Ol0O.addnsub_multiplier_pipeline_register1 = "UNREGISTERED",
		nl1Ol0O.addnsub_multiplier_pipeline_register3 = "UNREGISTERED",
		nl1Ol0O.addnsub_multiplier_register1 = "CLOCK0",
		nl1Ol0O.addnsub_multiplier_register3 = "CLOCK0",
		nl1Ol0O.chainout_aclr = "ACLR3",
		nl1Ol0O.chainout_adder = "NO",
		nl1Ol0O.chainout_register = "CLOCK0",
		nl1Ol0O.chainout_round_aclr = "ACLR3",
		nl1Ol0O.chainout_round_output_aclr = "ACLR3",
		nl1Ol0O.chainout_round_output_register = "CLOCK0",
		nl1Ol0O.chainout_round_pipeline_aclr = "ACLR3",
		nl1Ol0O.chainout_round_pipeline_register = "CLOCK0",
		nl1Ol0O.chainout_round_register = "CLOCK0",
		nl1Ol0O.chainout_rounding = "NO",
		nl1Ol0O.chainout_saturate_aclr = "ACLR3",
		nl1Ol0O.chainout_saturate_output_aclr = "ACLR3",
		nl1Ol0O.chainout_saturate_output_register = "CLOCK0",
		nl1Ol0O.chainout_saturate_pipeline_aclr = "ACLR3",
		nl1Ol0O.chainout_saturate_pipeline_register = "CLOCK0",
		nl1Ol0O.chainout_saturate_register = "CLOCK0",
		nl1Ol0O.chainout_saturation = "NO",
		nl1Ol0O.coef0_0 = 0,
		nl1Ol0O.coef0_1 = 0,
		nl1Ol0O.coef0_2 = 0,
		nl1Ol0O.coef0_3 = 0,
		nl1Ol0O.coef0_4 = 0,
		nl1Ol0O.coef0_5 = 0,
		nl1Ol0O.coef0_6 = 0,
		nl1Ol0O.coef0_7 = 0,
		nl1Ol0O.coef1_0 = 0,
		nl1Ol0O.coef1_1 = 0,
		nl1Ol0O.coef1_2 = 0,
		nl1Ol0O.coef1_3 = 0,
		nl1Ol0O.coef1_4 = 0,
		nl1Ol0O.coef1_5 = 0,
		nl1Ol0O.coef1_6 = 0,
		nl1Ol0O.coef1_7 = 0,
		nl1Ol0O.coef2_0 = 0,
		nl1Ol0O.coef2_1 = 0,
		nl1Ol0O.coef2_2 = 0,
		nl1Ol0O.coef2_3 = 0,
		nl1Ol0O.coef2_4 = 0,
		nl1Ol0O.coef2_5 = 0,
		nl1Ol0O.coef2_6 = 0,
		nl1Ol0O.coef2_7 = 0,
		nl1Ol0O.coef3_0 = 0,
		nl1Ol0O.coef3_1 = 0,
		nl1Ol0O.coef3_2 = 0,
		nl1Ol0O.coef3_3 = 0,
		nl1Ol0O.coef3_4 = 0,
		nl1Ol0O.coef3_5 = 0,
		nl1Ol0O.coef3_6 = 0,
		nl1Ol0O.coef3_7 = 0,
		nl1Ol0O.coefsel0_aclr = "ACLR0",
		nl1Ol0O.coefsel0_register = "CLOCK0",
		nl1Ol0O.coefsel1_aclr = "ACLR0",
		nl1Ol0O.coefsel1_register = "CLOCK0",
		nl1Ol0O.coefsel2_aclr = "ACLR0",
		nl1Ol0O.coefsel2_register = "CLOCK0",
		nl1Ol0O.coefsel3_aclr = "ACLR0",
		nl1Ol0O.coefsel3_register = "CLOCK0",
		nl1Ol0O.dsp_block_balancing = "AUTO",
		nl1Ol0O.extra_latency = 0,
		nl1Ol0O.input_aclr_a0 = "ACLR3",
		nl1Ol0O.input_aclr_a1 = "ACLR3",
		nl1Ol0O.input_aclr_a2 = "ACLR3",
		nl1Ol0O.input_aclr_a3 = "ACLR3",
		nl1Ol0O.input_aclr_b0 = "ACLR3",
		nl1Ol0O.input_aclr_b1 = "ACLR3",
		nl1Ol0O.input_aclr_b2 = "ACLR3",
		nl1Ol0O.input_aclr_b3 = "ACLR3",
		nl1Ol0O.input_aclr_c0 = "ACLR0",
		nl1Ol0O.input_register_a0 = "CLOCK0",
		nl1Ol0O.input_register_a1 = "CLOCK0",
		nl1Ol0O.input_register_a2 = "CLOCK0",
		nl1Ol0O.input_register_a3 = "CLOCK0",
		nl1Ol0O.input_register_b0 = "CLOCK0",
		nl1Ol0O.input_register_b1 = "CLOCK0",
		nl1Ol0O.input_register_b2 = "CLOCK0",
		nl1Ol0O.input_register_b3 = "CLOCK0",
		nl1Ol0O.input_register_c0 = "CLOCK0",
		nl1Ol0O.input_source_a0 = "DATAA",
		nl1Ol0O.input_source_a1 = "DATAA",
		nl1Ol0O.input_source_a2 = "DATAA",
		nl1Ol0O.input_source_a3 = "DATAA",
		nl1Ol0O.input_source_b0 = "DATAB",
		nl1Ol0O.input_source_b1 = "DATAB",
		nl1Ol0O.input_source_b2 = "DATAB",
		nl1Ol0O.input_source_b3 = "DATAB",
		nl1Ol0O.intended_device_family = "Cyclone III",
		nl1Ol0O.loadconst_value = 64,
		nl1Ol0O.mult01_round_aclr = "ACLR3",
		nl1Ol0O.mult01_round_register = "CLOCK0",
		nl1Ol0O.mult01_saturation_aclr = "ACLR2",
		nl1Ol0O.mult01_saturation_register = "CLOCK0",
		nl1Ol0O.mult23_round_aclr = "ACLR3",
		nl1Ol0O.mult23_round_register = "CLOCK0",
		nl1Ol0O.mult23_saturation_aclr = "ACLR3",
		nl1Ol0O.mult23_saturation_register = "CLOCK0",
		nl1Ol0O.multiplier01_rounding = "NO",
		nl1Ol0O.multiplier01_saturation = "NO",
		nl1Ol0O.multiplier1_direction = "ADD",
		nl1Ol0O.multiplier23_rounding = "NO",
		nl1Ol0O.multiplier23_saturation = "NO",
		nl1Ol0O.multiplier3_direction = "ADD",
		nl1Ol0O.multiplier_aclr0 = "ACLR3",
		nl1Ol0O.multiplier_aclr1 = "ACLR3",
		nl1Ol0O.multiplier_aclr2 = "ACLR3",
		nl1Ol0O.multiplier_aclr3 = "ACLR3",
		nl1Ol0O.multiplier_register0 = "CLOCK0",
		nl1Ol0O.multiplier_register1 = "CLOCK0",
		nl1Ol0O.multiplier_register2 = "CLOCK0",
		nl1Ol0O.multiplier_register3 = "CLOCK0",
		nl1Ol0O.number_of_multipliers = 1,
		nl1Ol0O.output_aclr = "ACLR0",
		nl1Ol0O.output_register = "CLOCK0",
		nl1Ol0O.output_round_aclr = "ACLR3",
		nl1Ol0O.output_round_pipeline_aclr = "ACLR3",
		nl1Ol0O.output_round_pipeline_register = "CLOCK0",
		nl1Ol0O.output_round_register = "CLOCK0",
		nl1Ol0O.output_round_type = "NEAREST_INTEGER",
		nl1Ol0O.output_rounding = "NO",
		nl1Ol0O.output_saturate_aclr = "ACLR3",
		nl1Ol0O.output_saturate_pipeline_aclr = "ACLR3",
		nl1Ol0O.output_saturate_pipeline_register = "CLOCK0",
		nl1Ol0O.output_saturate_register = "CLOCK0",
		nl1Ol0O.output_saturate_type = "ASYMMETRIC",
		nl1Ol0O.output_saturation = "NO",
		nl1Ol0O.port_addnsub1 = "PORT_UNUSED",
		nl1Ol0O.port_addnsub3 = "PORT_UNUSED",
		nl1Ol0O.port_chainout_sat_is_overflow = "PORT_UNUSED",
		nl1Ol0O.port_output_is_overflow = "PORT_UNUSED",
		nl1Ol0O.port_signa = "PORT_CONNECTIVITY",
		nl1Ol0O.port_signb = "PORT_CONNECTIVITY",
		nl1Ol0O.preadder_direction_0 = "ADD",
		nl1Ol0O.preadder_direction_1 = "ADD",
		nl1Ol0O.preadder_direction_2 = "ADD",
		nl1Ol0O.preadder_direction_3 = "ADD",
		nl1Ol0O.preadder_mode = "SIMPLE",
		nl1Ol0O.representation_a = "UNSIGNED",
		nl1Ol0O.representation_b = "UNSIGNED",
		nl1Ol0O.rotate_aclr = "ACLR3",
		nl1Ol0O.rotate_output_aclr = "ACLR3",
		nl1Ol0O.rotate_output_register = "CLOCK0",
		nl1Ol0O.rotate_pipeline_aclr = "ACLR3",
		nl1Ol0O.rotate_pipeline_register = "CLOCK0",
		nl1Ol0O.rotate_register = "CLOCK0",
		nl1Ol0O.scanouta_aclr = "ACLR3",
		nl1Ol0O.scanouta_register = "UNREGISTERED",
		nl1Ol0O.shift_mode = "NO",
		nl1Ol0O.shift_right_aclr = "ACLR3",
		nl1Ol0O.shift_right_output_aclr = "ACLR3",
		nl1Ol0O.shift_right_output_register = "CLOCK0",
		nl1Ol0O.shift_right_pipeline_aclr = "ACLR3",
		nl1Ol0O.shift_right_pipeline_register = "CLOCK0",
		nl1Ol0O.shift_right_register = "CLOCK0",
		nl1Ol0O.signed_aclr_a = "ACLR3",
		nl1Ol0O.signed_aclr_b = "ACLR3",
		nl1Ol0O.signed_pipeline_aclr_a = "ACLR3",
		nl1Ol0O.signed_pipeline_aclr_b = "ACLR3",
		nl1Ol0O.signed_pipeline_register_a = "UNREGISTERED",
		nl1Ol0O.signed_pipeline_register_b = "UNREGISTERED",
		nl1Ol0O.signed_register_a = "CLOCK0",
		nl1Ol0O.signed_register_b = "CLOCK0",
		nl1Ol0O.systolic_aclr1 = "ACLR0",
		nl1Ol0O.systolic_aclr3 = "ACLR0",
		nl1Ol0O.systolic_delay1 = "UNREGISTERED",
		nl1Ol0O.systolic_delay3 = "UNREGISTERED",
		nl1Ol0O.width_a = 9,
		nl1Ol0O.width_b = 9,
		nl1Ol0O.width_c = 22,
		nl1Ol0O.width_chainin = 1,
		nl1Ol0O.width_coef = 18,
		nl1Ol0O.width_msb = 17,
		nl1Ol0O.width_result = 18,
		nl1Ol0O.width_saturate_sign = 1,
		nl1Ol0O.zero_chainout_output_aclr = "ACLR3",
		nl1Ol0O.zero_chainout_output_register = "CLOCK0",
		nl1Ol0O.zero_loopback_aclr = "ACLR3",
		nl1Ol0O.zero_loopback_output_aclr = "ACLR3",
		nl1Ol0O.zero_loopback_output_register = "CLOCK0",
		nl1Ol0O.zero_loopback_pipeline_aclr = "ACLR3",
		nl1Ol0O.zero_loopback_pipeline_register = "CLOCK0",
		nl1Ol0O.zero_loopback_register = "CLOCK0";
	altmult_add   nl1OllO
	( 
	.chainout_sat_overflow(),
	.clock0(clock),
	.dataa({nl1O00i, nl1O01O, nl1O01l, nl1O01i, nl1O1OO, nl1O1Ol, nl1O1Oi, nl1O1lO, nl1O00O}),
	.datab({1'b0, nli000l, nli001O, nli001l, nli001i, nli01OO, nli01Ol, nli01Oi, nli01lO}),
	.ena0(((~ ni1iili) & ((n010l | nl1OO1l) | nl1OlOi))),
	.mult0_is_saturated(),
	.mult1_is_saturated(),
	.mult2_is_saturated(),
	.mult3_is_saturated(),
	.overflow(),
	.result(wire_nl1OllO_result),
	.scanouta(),
	.scanoutb(),
	.signa(1'b0),
	.signb(1'b0),
	.accum_sload(),
	.aclr0(),
	.aclr1(),
	.aclr2(),
	.aclr3(),
	.addnsub1(),
	.addnsub1_round(),
	.addnsub3(),
	.addnsub3_round(),
	.chainin(),
	.chainout_round(),
	.chainout_saturate(),
	.clock1(),
	.clock2(),
	.clock3(),
	.coefsel0(),
	.coefsel1(),
	.coefsel2(),
	.coefsel3(),
	.datac(),
	.ena1(),
	.ena2(),
	.ena3(),
	.mult01_round(),
	.mult01_saturation(),
	.mult23_round(),
	.mult23_saturation(),
	.output_round(),
	.output_saturate(),
	.rotate(),
	.scanina(),
	.scaninb(),
	.shift_right(),
	.sourcea(),
	.sourceb(),
	.zero_chainout(),
	.zero_loopback()
	);
	defparam
		nl1OllO.accum_direction = "ADD",
		nl1OllO.accum_sload_aclr = "ACLR3",
		nl1OllO.accum_sload_pipeline_aclr = "ACLR3",
		nl1OllO.accum_sload_pipeline_register = "CLOCK0",
		nl1OllO.accum_sload_register = "CLOCK0",
		nl1OllO.accumulator = "NO",
		nl1OllO.adder1_rounding = "NO",
		nl1OllO.adder3_rounding = "NO",
		nl1OllO.addnsub1_round_aclr = "ACLR3",
		nl1OllO.addnsub1_round_pipeline_aclr = "ACLR3",
		nl1OllO.addnsub1_round_pipeline_register = "CLOCK0",
		nl1OllO.addnsub1_round_register = "CLOCK0",
		nl1OllO.addnsub3_round_aclr = "ACLR3",
		nl1OllO.addnsub3_round_pipeline_aclr = "ACLR3",
		nl1OllO.addnsub3_round_pipeline_register = "CLOCK0",
		nl1OllO.addnsub3_round_register = "CLOCK0",
		nl1OllO.addnsub_multiplier_aclr1 = "ACLR3",
		nl1OllO.addnsub_multiplier_aclr3 = "ACLR3",
		nl1OllO.addnsub_multiplier_pipeline_aclr1 = "ACLR3",
		nl1OllO.addnsub_multiplier_pipeline_aclr3 = "ACLR3",
		nl1OllO.addnsub_multiplier_pipeline_register1 = "UNREGISTERED",
		nl1OllO.addnsub_multiplier_pipeline_register3 = "UNREGISTERED",
		nl1OllO.addnsub_multiplier_register1 = "CLOCK0",
		nl1OllO.addnsub_multiplier_register3 = "CLOCK0",
		nl1OllO.chainout_aclr = "ACLR3",
		nl1OllO.chainout_adder = "NO",
		nl1OllO.chainout_register = "CLOCK0",
		nl1OllO.chainout_round_aclr = "ACLR3",
		nl1OllO.chainout_round_output_aclr = "ACLR3",
		nl1OllO.chainout_round_output_register = "CLOCK0",
		nl1OllO.chainout_round_pipeline_aclr = "ACLR3",
		nl1OllO.chainout_round_pipeline_register = "CLOCK0",
		nl1OllO.chainout_round_register = "CLOCK0",
		nl1OllO.chainout_rounding = "NO",
		nl1OllO.chainout_saturate_aclr = "ACLR3",
		nl1OllO.chainout_saturate_output_aclr = "ACLR3",
		nl1OllO.chainout_saturate_output_register = "CLOCK0",
		nl1OllO.chainout_saturate_pipeline_aclr = "ACLR3",
		nl1OllO.chainout_saturate_pipeline_register = "CLOCK0",
		nl1OllO.chainout_saturate_register = "CLOCK0",
		nl1OllO.chainout_saturation = "NO",
		nl1OllO.coef0_0 = 0,
		nl1OllO.coef0_1 = 0,
		nl1OllO.coef0_2 = 0,
		nl1OllO.coef0_3 = 0,
		nl1OllO.coef0_4 = 0,
		nl1OllO.coef0_5 = 0,
		nl1OllO.coef0_6 = 0,
		nl1OllO.coef0_7 = 0,
		nl1OllO.coef1_0 = 0,
		nl1OllO.coef1_1 = 0,
		nl1OllO.coef1_2 = 0,
		nl1OllO.coef1_3 = 0,
		nl1OllO.coef1_4 = 0,
		nl1OllO.coef1_5 = 0,
		nl1OllO.coef1_6 = 0,
		nl1OllO.coef1_7 = 0,
		nl1OllO.coef2_0 = 0,
		nl1OllO.coef2_1 = 0,
		nl1OllO.coef2_2 = 0,
		nl1OllO.coef2_3 = 0,
		nl1OllO.coef2_4 = 0,
		nl1OllO.coef2_5 = 0,
		nl1OllO.coef2_6 = 0,
		nl1OllO.coef2_7 = 0,
		nl1OllO.coef3_0 = 0,
		nl1OllO.coef3_1 = 0,
		nl1OllO.coef3_2 = 0,
		nl1OllO.coef3_3 = 0,
		nl1OllO.coef3_4 = 0,
		nl1OllO.coef3_5 = 0,
		nl1OllO.coef3_6 = 0,
		nl1OllO.coef3_7 = 0,
		nl1OllO.coefsel0_aclr = "ACLR0",
		nl1OllO.coefsel0_register = "CLOCK0",
		nl1OllO.coefsel1_aclr = "ACLR0",
		nl1OllO.coefsel1_register = "CLOCK0",
		nl1OllO.coefsel2_aclr = "ACLR0",
		nl1OllO.coefsel2_register = "CLOCK0",
		nl1OllO.coefsel3_aclr = "ACLR0",
		nl1OllO.coefsel3_register = "CLOCK0",
		nl1OllO.dsp_block_balancing = "AUTO",
		nl1OllO.extra_latency = 0,
		nl1OllO.input_aclr_a0 = "ACLR3",
		nl1OllO.input_aclr_a1 = "ACLR3",
		nl1OllO.input_aclr_a2 = "ACLR3",
		nl1OllO.input_aclr_a3 = "ACLR3",
		nl1OllO.input_aclr_b0 = "ACLR3",
		nl1OllO.input_aclr_b1 = "ACLR3",
		nl1OllO.input_aclr_b2 = "ACLR3",
		nl1OllO.input_aclr_b3 = "ACLR3",
		nl1OllO.input_aclr_c0 = "ACLR0",
		nl1OllO.input_register_a0 = "CLOCK0",
		nl1OllO.input_register_a1 = "CLOCK0",
		nl1OllO.input_register_a2 = "CLOCK0",
		nl1OllO.input_register_a3 = "CLOCK0",
		nl1OllO.input_register_b0 = "CLOCK0",
		nl1OllO.input_register_b1 = "CLOCK0",
		nl1OllO.input_register_b2 = "CLOCK0",
		nl1OllO.input_register_b3 = "CLOCK0",
		nl1OllO.input_register_c0 = "CLOCK0",
		nl1OllO.input_source_a0 = "DATAA",
		nl1OllO.input_source_a1 = "DATAA",
		nl1OllO.input_source_a2 = "DATAA",
		nl1OllO.input_source_a3 = "DATAA",
		nl1OllO.input_source_b0 = "DATAB",
		nl1OllO.input_source_b1 = "DATAB",
		nl1OllO.input_source_b2 = "DATAB",
		nl1OllO.input_source_b3 = "DATAB",
		nl1OllO.intended_device_family = "Cyclone III",
		nl1OllO.loadconst_value = 64,
		nl1OllO.mult01_round_aclr = "ACLR3",
		nl1OllO.mult01_round_register = "CLOCK0",
		nl1OllO.mult01_saturation_aclr = "ACLR2",
		nl1OllO.mult01_saturation_register = "CLOCK0",
		nl1OllO.mult23_round_aclr = "ACLR3",
		nl1OllO.mult23_round_register = "CLOCK0",
		nl1OllO.mult23_saturation_aclr = "ACLR3",
		nl1OllO.mult23_saturation_register = "CLOCK0",
		nl1OllO.multiplier01_rounding = "NO",
		nl1OllO.multiplier01_saturation = "NO",
		nl1OllO.multiplier1_direction = "ADD",
		nl1OllO.multiplier23_rounding = "NO",
		nl1OllO.multiplier23_saturation = "NO",
		nl1OllO.multiplier3_direction = "ADD",
		nl1OllO.multiplier_aclr0 = "ACLR3",
		nl1OllO.multiplier_aclr1 = "ACLR3",
		nl1OllO.multiplier_aclr2 = "ACLR3",
		nl1OllO.multiplier_aclr3 = "ACLR3",
		nl1OllO.multiplier_register0 = "CLOCK0",
		nl1OllO.multiplier_register1 = "CLOCK0",
		nl1OllO.multiplier_register2 = "CLOCK0",
		nl1OllO.multiplier_register3 = "CLOCK0",
		nl1OllO.number_of_multipliers = 1,
		nl1OllO.output_aclr = "ACLR0",
		nl1OllO.output_register = "CLOCK0",
		nl1OllO.output_round_aclr = "ACLR3",
		nl1OllO.output_round_pipeline_aclr = "ACLR3",
		nl1OllO.output_round_pipeline_register = "CLOCK0",
		nl1OllO.output_round_register = "CLOCK0",
		nl1OllO.output_round_type = "NEAREST_INTEGER",
		nl1OllO.output_rounding = "NO",
		nl1OllO.output_saturate_aclr = "ACLR3",
		nl1OllO.output_saturate_pipeline_aclr = "ACLR3",
		nl1OllO.output_saturate_pipeline_register = "CLOCK0",
		nl1OllO.output_saturate_register = "CLOCK0",
		nl1OllO.output_saturate_type = "ASYMMETRIC",
		nl1OllO.output_saturation = "NO",
		nl1OllO.port_addnsub1 = "PORT_UNUSED",
		nl1OllO.port_addnsub3 = "PORT_UNUSED",
		nl1OllO.port_chainout_sat_is_overflow = "PORT_UNUSED",
		nl1OllO.port_output_is_overflow = "PORT_UNUSED",
		nl1OllO.port_signa = "PORT_CONNECTIVITY",
		nl1OllO.port_signb = "PORT_CONNECTIVITY",
		nl1OllO.preadder_direction_0 = "ADD",
		nl1OllO.preadder_direction_1 = "ADD",
		nl1OllO.preadder_direction_2 = "ADD",
		nl1OllO.preadder_direction_3 = "ADD",
		nl1OllO.preadder_mode = "SIMPLE",
		nl1OllO.representation_a = "UNSIGNED",
		nl1OllO.representation_b = "UNSIGNED",
		nl1OllO.rotate_aclr = "ACLR3",
		nl1OllO.rotate_output_aclr = "ACLR3",
		nl1OllO.rotate_output_register = "CLOCK0",
		nl1OllO.rotate_pipeline_aclr = "ACLR3",
		nl1OllO.rotate_pipeline_register = "CLOCK0",
		nl1OllO.rotate_register = "CLOCK0",
		nl1OllO.scanouta_aclr = "ACLR3",
		nl1OllO.scanouta_register = "UNREGISTERED",
		nl1OllO.shift_mode = "NO",
		nl1OllO.shift_right_aclr = "ACLR3",
		nl1OllO.shift_right_output_aclr = "ACLR3",
		nl1OllO.shift_right_output_register = "CLOCK0",
		nl1OllO.shift_right_pipeline_aclr = "ACLR3",
		nl1OllO.shift_right_pipeline_register = "CLOCK0",
		nl1OllO.shift_right_register = "CLOCK0",
		nl1OllO.signed_aclr_a = "ACLR3",
		nl1OllO.signed_aclr_b = "ACLR3",
		nl1OllO.signed_pipeline_aclr_a = "ACLR3",
		nl1OllO.signed_pipeline_aclr_b = "ACLR3",
		nl1OllO.signed_pipeline_register_a = "UNREGISTERED",
		nl1OllO.signed_pipeline_register_b = "UNREGISTERED",
		nl1OllO.signed_register_a = "CLOCK0",
		nl1OllO.signed_register_b = "CLOCK0",
		nl1OllO.systolic_aclr1 = "ACLR0",
		nl1OllO.systolic_aclr3 = "ACLR0",
		nl1OllO.systolic_delay1 = "UNREGISTERED",
		nl1OllO.systolic_delay3 = "UNREGISTERED",
		nl1OllO.width_a = 9,
		nl1OllO.width_b = 9,
		nl1OllO.width_c = 22,
		nl1OllO.width_chainin = 1,
		nl1OllO.width_coef = 18,
		nl1OllO.width_msb = 17,
		nl1OllO.width_result = 18,
		nl1OllO.width_saturate_sign = 1,
		nl1OllO.zero_chainout_output_aclr = "ACLR3",
		nl1OllO.zero_chainout_output_register = "CLOCK0",
		nl1OllO.zero_loopback_aclr = "ACLR3",
		nl1OllO.zero_loopback_output_aclr = "ACLR3",
		nl1OllO.zero_loopback_output_register = "CLOCK0",
		nl1OllO.zero_loopback_pipeline_aclr = "ACLR3",
		nl1OllO.zero_loopback_pipeline_register = "CLOCK0",
		nl1OllO.zero_loopback_register = "CLOCK0";
	altmult_add   nl1OO1O
	( 
	.chainout_sat_overflow(),
	.clock0(clock),
	.dataa({nl1O00i, nl1O01O, nl1O01l, nl1O01i, nl1O1OO, nl1O1Ol, nl1O1Oi, nl1O1lO, nl1O00O}),
	.datab({1'b0, nli01li, nli01il, nli01ii, nli010O, nli010l, nli010i, nli011O, nli011l}),
	.ena0(((~ ni1iili) & ((n010l | nl1OOiO) | nl1OO0i))),
	.mult0_is_saturated(),
	.mult1_is_saturated(),
	.mult2_is_saturated(),
	.mult3_is_saturated(),
	.overflow(),
	.result(wire_nl1OO1O_result),
	.scanouta(),
	.scanoutb(),
	.signa(1'b0),
	.signb(1'b0),
	.accum_sload(),
	.aclr0(),
	.aclr1(),
	.aclr2(),
	.aclr3(),
	.addnsub1(),
	.addnsub1_round(),
	.addnsub3(),
	.addnsub3_round(),
	.chainin(),
	.chainout_round(),
	.chainout_saturate(),
	.clock1(),
	.clock2(),
	.clock3(),
	.coefsel0(),
	.coefsel1(),
	.coefsel2(),
	.coefsel3(),
	.datac(),
	.ena1(),
	.ena2(),
	.ena3(),
	.mult01_round(),
	.mult01_saturation(),
	.mult23_round(),
	.mult23_saturation(),
	.output_round(),
	.output_saturate(),
	.rotate(),
	.scanina(),
	.scaninb(),
	.shift_right(),
	.sourcea(),
	.sourceb(),
	.zero_chainout(),
	.zero_loopback()
	);
	defparam
		nl1OO1O.accum_direction = "ADD",
		nl1OO1O.accum_sload_aclr = "ACLR3",
		nl1OO1O.accum_sload_pipeline_aclr = "ACLR3",
		nl1OO1O.accum_sload_pipeline_register = "CLOCK0",
		nl1OO1O.accum_sload_register = "CLOCK0",
		nl1OO1O.accumulator = "NO",
		nl1OO1O.adder1_rounding = "NO",
		nl1OO1O.adder3_rounding = "NO",
		nl1OO1O.addnsub1_round_aclr = "ACLR3",
		nl1OO1O.addnsub1_round_pipeline_aclr = "ACLR3",
		nl1OO1O.addnsub1_round_pipeline_register = "CLOCK0",
		nl1OO1O.addnsub1_round_register = "CLOCK0",
		nl1OO1O.addnsub3_round_aclr = "ACLR3",
		nl1OO1O.addnsub3_round_pipeline_aclr = "ACLR3",
		nl1OO1O.addnsub3_round_pipeline_register = "CLOCK0",
		nl1OO1O.addnsub3_round_register = "CLOCK0",
		nl1OO1O.addnsub_multiplier_aclr1 = "ACLR3",
		nl1OO1O.addnsub_multiplier_aclr3 = "ACLR3",
		nl1OO1O.addnsub_multiplier_pipeline_aclr1 = "ACLR3",
		nl1OO1O.addnsub_multiplier_pipeline_aclr3 = "ACLR3",
		nl1OO1O.addnsub_multiplier_pipeline_register1 = "UNREGISTERED",
		nl1OO1O.addnsub_multiplier_pipeline_register3 = "UNREGISTERED",
		nl1OO1O.addnsub_multiplier_register1 = "CLOCK0",
		nl1OO1O.addnsub_multiplier_register3 = "CLOCK0",
		nl1OO1O.chainout_aclr = "ACLR3",
		nl1OO1O.chainout_adder = "NO",
		nl1OO1O.chainout_register = "CLOCK0",
		nl1OO1O.chainout_round_aclr = "ACLR3",
		nl1OO1O.chainout_round_output_aclr = "ACLR3",
		nl1OO1O.chainout_round_output_register = "CLOCK0",
		nl1OO1O.chainout_round_pipeline_aclr = "ACLR3",
		nl1OO1O.chainout_round_pipeline_register = "CLOCK0",
		nl1OO1O.chainout_round_register = "CLOCK0",
		nl1OO1O.chainout_rounding = "NO",
		nl1OO1O.chainout_saturate_aclr = "ACLR3",
		nl1OO1O.chainout_saturate_output_aclr = "ACLR3",
		nl1OO1O.chainout_saturate_output_register = "CLOCK0",
		nl1OO1O.chainout_saturate_pipeline_aclr = "ACLR3",
		nl1OO1O.chainout_saturate_pipeline_register = "CLOCK0",
		nl1OO1O.chainout_saturate_register = "CLOCK0",
		nl1OO1O.chainout_saturation = "NO",
		nl1OO1O.coef0_0 = 0,
		nl1OO1O.coef0_1 = 0,
		nl1OO1O.coef0_2 = 0,
		nl1OO1O.coef0_3 = 0,
		nl1OO1O.coef0_4 = 0,
		nl1OO1O.coef0_5 = 0,
		nl1OO1O.coef0_6 = 0,
		nl1OO1O.coef0_7 = 0,
		nl1OO1O.coef1_0 = 0,
		nl1OO1O.coef1_1 = 0,
		nl1OO1O.coef1_2 = 0,
		nl1OO1O.coef1_3 = 0,
		nl1OO1O.coef1_4 = 0,
		nl1OO1O.coef1_5 = 0,
		nl1OO1O.coef1_6 = 0,
		nl1OO1O.coef1_7 = 0,
		nl1OO1O.coef2_0 = 0,
		nl1OO1O.coef2_1 = 0,
		nl1OO1O.coef2_2 = 0,
		nl1OO1O.coef2_3 = 0,
		nl1OO1O.coef2_4 = 0,
		nl1OO1O.coef2_5 = 0,
		nl1OO1O.coef2_6 = 0,
		nl1OO1O.coef2_7 = 0,
		nl1OO1O.coef3_0 = 0,
		nl1OO1O.coef3_1 = 0,
		nl1OO1O.coef3_2 = 0,
		nl1OO1O.coef3_3 = 0,
		nl1OO1O.coef3_4 = 0,
		nl1OO1O.coef3_5 = 0,
		nl1OO1O.coef3_6 = 0,
		nl1OO1O.coef3_7 = 0,
		nl1OO1O.coefsel0_aclr = "ACLR0",
		nl1OO1O.coefsel0_register = "CLOCK0",
		nl1OO1O.coefsel1_aclr = "ACLR0",
		nl1OO1O.coefsel1_register = "CLOCK0",
		nl1OO1O.coefsel2_aclr = "ACLR0",
		nl1OO1O.coefsel2_register = "CLOCK0",
		nl1OO1O.coefsel3_aclr = "ACLR0",
		nl1OO1O.coefsel3_register = "CLOCK0",
		nl1OO1O.dsp_block_balancing = "AUTO",
		nl1OO1O.extra_latency = 0,
		nl1OO1O.input_aclr_a0 = "ACLR3",
		nl1OO1O.input_aclr_a1 = "ACLR3",
		nl1OO1O.input_aclr_a2 = "ACLR3",
		nl1OO1O.input_aclr_a3 = "ACLR3",
		nl1OO1O.input_aclr_b0 = "ACLR3",
		nl1OO1O.input_aclr_b1 = "ACLR3",
		nl1OO1O.input_aclr_b2 = "ACLR3",
		nl1OO1O.input_aclr_b3 = "ACLR3",
		nl1OO1O.input_aclr_c0 = "ACLR0",
		nl1OO1O.input_register_a0 = "CLOCK0",
		nl1OO1O.input_register_a1 = "CLOCK0",
		nl1OO1O.input_register_a2 = "CLOCK0",
		nl1OO1O.input_register_a3 = "CLOCK0",
		nl1OO1O.input_register_b0 = "CLOCK0",
		nl1OO1O.input_register_b1 = "CLOCK0",
		nl1OO1O.input_register_b2 = "CLOCK0",
		nl1OO1O.input_register_b3 = "CLOCK0",
		nl1OO1O.input_register_c0 = "CLOCK0",
		nl1OO1O.input_source_a0 = "DATAA",
		nl1OO1O.input_source_a1 = "DATAA",
		nl1OO1O.input_source_a2 = "DATAA",
		nl1OO1O.input_source_a3 = "DATAA",
		nl1OO1O.input_source_b0 = "DATAB",
		nl1OO1O.input_source_b1 = "DATAB",
		nl1OO1O.input_source_b2 = "DATAB",
		nl1OO1O.input_source_b3 = "DATAB",
		nl1OO1O.intended_device_family = "Cyclone III",
		nl1OO1O.loadconst_value = 64,
		nl1OO1O.mult01_round_aclr = "ACLR3",
		nl1OO1O.mult01_round_register = "CLOCK0",
		nl1OO1O.mult01_saturation_aclr = "ACLR2",
		nl1OO1O.mult01_saturation_register = "CLOCK0",
		nl1OO1O.mult23_round_aclr = "ACLR3",
		nl1OO1O.mult23_round_register = "CLOCK0",
		nl1OO1O.mult23_saturation_aclr = "ACLR3",
		nl1OO1O.mult23_saturation_register = "CLOCK0",
		nl1OO1O.multiplier01_rounding = "NO",
		nl1OO1O.multiplier01_saturation = "NO",
		nl1OO1O.multiplier1_direction = "ADD",
		nl1OO1O.multiplier23_rounding = "NO",
		nl1OO1O.multiplier23_saturation = "NO",
		nl1OO1O.multiplier3_direction = "ADD",
		nl1OO1O.multiplier_aclr0 = "ACLR3",
		nl1OO1O.multiplier_aclr1 = "ACLR3",
		nl1OO1O.multiplier_aclr2 = "ACLR3",
		nl1OO1O.multiplier_aclr3 = "ACLR3",
		nl1OO1O.multiplier_register0 = "CLOCK0",
		nl1OO1O.multiplier_register1 = "CLOCK0",
		nl1OO1O.multiplier_register2 = "CLOCK0",
		nl1OO1O.multiplier_register3 = "CLOCK0",
		nl1OO1O.number_of_multipliers = 1,
		nl1OO1O.output_aclr = "ACLR0",
		nl1OO1O.output_register = "CLOCK0",
		nl1OO1O.output_round_aclr = "ACLR3",
		nl1OO1O.output_round_pipeline_aclr = "ACLR3",
		nl1OO1O.output_round_pipeline_register = "CLOCK0",
		nl1OO1O.output_round_register = "CLOCK0",
		nl1OO1O.output_round_type = "NEAREST_INTEGER",
		nl1OO1O.output_rounding = "NO",
		nl1OO1O.output_saturate_aclr = "ACLR3",
		nl1OO1O.output_saturate_pipeline_aclr = "ACLR3",
		nl1OO1O.output_saturate_pipeline_register = "CLOCK0",
		nl1OO1O.output_saturate_register = "CLOCK0",
		nl1OO1O.output_saturate_type = "ASYMMETRIC",
		nl1OO1O.output_saturation = "NO",
		nl1OO1O.port_addnsub1 = "PORT_UNUSED",
		nl1OO1O.port_addnsub3 = "PORT_UNUSED",
		nl1OO1O.port_chainout_sat_is_overflow = "PORT_UNUSED",
		nl1OO1O.port_output_is_overflow = "PORT_UNUSED",
		nl1OO1O.port_signa = "PORT_CONNECTIVITY",
		nl1OO1O.port_signb = "PORT_CONNECTIVITY",
		nl1OO1O.preadder_direction_0 = "ADD",
		nl1OO1O.preadder_direction_1 = "ADD",
		nl1OO1O.preadder_direction_2 = "ADD",
		nl1OO1O.preadder_direction_3 = "ADD",
		nl1OO1O.preadder_mode = "SIMPLE",
		nl1OO1O.representation_a = "UNSIGNED",
		nl1OO1O.representation_b = "UNSIGNED",
		nl1OO1O.rotate_aclr = "ACLR3",
		nl1OO1O.rotate_output_aclr = "ACLR3",
		nl1OO1O.rotate_output_register = "CLOCK0",
		nl1OO1O.rotate_pipeline_aclr = "ACLR3",
		nl1OO1O.rotate_pipeline_register = "CLOCK0",
		nl1OO1O.rotate_register = "CLOCK0",
		nl1OO1O.scanouta_aclr = "ACLR3",
		nl1OO1O.scanouta_register = "UNREGISTERED",
		nl1OO1O.shift_mode = "NO",
		nl1OO1O.shift_right_aclr = "ACLR3",
		nl1OO1O.shift_right_output_aclr = "ACLR3",
		nl1OO1O.shift_right_output_register = "CLOCK0",
		nl1OO1O.shift_right_pipeline_aclr = "ACLR3",
		nl1OO1O.shift_right_pipeline_register = "CLOCK0",
		nl1OO1O.shift_right_register = "CLOCK0",
		nl1OO1O.signed_aclr_a = "ACLR3",
		nl1OO1O.signed_aclr_b = "ACLR3",
		nl1OO1O.signed_pipeline_aclr_a = "ACLR3",
		nl1OO1O.signed_pipeline_aclr_b = "ACLR3",
		nl1OO1O.signed_pipeline_register_a = "UNREGISTERED",
		nl1OO1O.signed_pipeline_register_b = "UNREGISTERED",
		nl1OO1O.signed_register_a = "CLOCK0",
		nl1OO1O.signed_register_b = "CLOCK0",
		nl1OO1O.systolic_aclr1 = "ACLR0",
		nl1OO1O.systolic_aclr3 = "ACLR0",
		nl1OO1O.systolic_delay1 = "UNREGISTERED",
		nl1OO1O.systolic_delay3 = "UNREGISTERED",
		nl1OO1O.width_a = 9,
		nl1OO1O.width_b = 9,
		nl1OO1O.width_c = 22,
		nl1OO1O.width_chainin = 1,
		nl1OO1O.width_coef = 18,
		nl1OO1O.width_msb = 17,
		nl1OO1O.width_result = 18,
		nl1OO1O.width_saturate_sign = 1,
		nl1OO1O.zero_chainout_output_aclr = "ACLR3",
		nl1OO1O.zero_chainout_output_register = "CLOCK0",
		nl1OO1O.zero_loopback_aclr = "ACLR3",
		nl1OO1O.zero_loopback_output_aclr = "ACLR3",
		nl1OO1O.zero_loopback_output_register = "CLOCK0",
		nl1OO1O.zero_loopback_pipeline_aclr = "ACLR3",
		nl1OO1O.zero_loopback_pipeline_register = "CLOCK0",
		nl1OO1O.zero_loopback_register = "CLOCK0";
	altsyncram   niOl0il
	( 
	.address_a({wire_niOl1li_dataout, wire_niOl1iO_dataout, wire_niOl1il_dataout, wire_niOl1ii_dataout, wire_niOl10O_dataout, wire_niOl10l_dataout}),
	.address_b({control_av_address[5:0]}),
	.clock0(clock),
	.clock1(clock),
	.clocken0(ni11Oll),
	.clocken1(1'b1),
	.data_a({{15{1'b0}}, n0O0O}),
	.data_b({control_av_writedata[15:0]}),
	.eccstatus(),
	.q_a(wire_niOl0il_q_a),
	.q_b(wire_niOl0il_q_b),
	.wren_a((n0Oii & n0O0l)),
	.wren_b((control_av_chipselect & control_av_write)),
	.aclr0(),
	.aclr1(),
	.addressstall_a(),
	.addressstall_b(),
	.byteena_a(),
	.byteena_b(),
	.clocken2(),
	.clocken3(),
	.rden_a(),
	.rden_b()
	);
	defparam
		niOl0il.address_aclr_a = "NONE",
		niOl0il.address_aclr_b = "NONE",
		niOl0il.address_reg_b = "CLOCK1",
		niOl0il.byte_size = 8,
		niOl0il.byteena_aclr_a = "NONE",
		niOl0il.byteena_aclr_b = "NONE",
		niOl0il.byteena_reg_b = "CLOCK1",
		niOl0il.clock_enable_core_a = "USE_INPUT_CLKEN",
		niOl0il.clock_enable_core_b = "USE_INPUT_CLKEN",
		niOl0il.clock_enable_input_a = "NORMAL",
		niOl0il.clock_enable_input_b = "NORMAL",
		niOl0il.clock_enable_output_a = "NORMAL",
		niOl0il.clock_enable_output_b = "NORMAL",
		niOl0il.ecc_pipeline_stage_enabled = "FALSE",
		niOl0il.enable_ecc = "FALSE",
		niOl0il.indata_aclr_a = "NONE",
		niOl0il.indata_aclr_b = "NONE",
		niOl0il.indata_reg_b = "CLOCK1",
		niOl0il.init_file = "UNUSED",
		niOl0il.init_file_layout = "PORT_A",
		niOl0il.intended_device_family = "Cyclone III",
		niOl0il.numwords_a = 47,
		niOl0il.numwords_b = 47,
		niOl0il.operation_mode = "BIDIR_DUAL_PORT",
		niOl0il.outdata_aclr_a = "NONE",
		niOl0il.outdata_aclr_b = "NONE",
		niOl0il.outdata_reg_a = "CLOCK0",
		niOl0il.outdata_reg_b = "CLOCK1",
		niOl0il.ram_block_type = "AUTO",
		niOl0il.rdcontrol_aclr_b = "NONE",
		niOl0il.rdcontrol_reg_b = "CLOCK1",
		niOl0il.read_during_write_mode_mixed_ports = "DONT_CARE",
		niOl0il.read_during_write_mode_port_a = "NEW_DATA_NO_NBE_READ",
		niOl0il.read_during_write_mode_port_b = "NEW_DATA_NO_NBE_READ",
		niOl0il.width_a = 16,
		niOl0il.width_b = 16,
		niOl0il.width_byteena_a = 1,
		niOl0il.width_byteena_b = 1,
		niOl0il.width_eccstatus = 3,
		niOl0il.widthad_a = 6,
		niOl0il.widthad_b = 6,
		niOl0il.wrcontrol_aclr_a = "NONE",
		niOl0il.wrcontrol_aclr_b = "NONE",
		niOl0il.wrcontrol_wraddress_reg_b = "CLOCK1",
		niOl0il.lpm_hint = "WIDTH_BYTEENA=1";
	initial
		ni1i00l63 = 0;
	always @ ( posedge clock)
		  ni1i00l63 <= ni1i00l64;
	event ni1i00l63_event;
	initial
		#1 ->ni1i00l63_event;
	always @(ni1i00l63_event)
		ni1i00l63 <= {1{1'b1}};
	initial
		ni1i00l64 = 0;
	always @ ( posedge clock)
		  ni1i00l64 <= ni1i00l63;
	initial
		ni1i00O61 = 0;
	always @ ( posedge clock)
		  ni1i00O61 <= ni1i00O62;
	event ni1i00O61_event;
	initial
		#1 ->ni1i00O61_event;
	always @(ni1i00O61_event)
		ni1i00O61 <= {1{1'b1}};
	initial
		ni1i00O62 = 0;
	always @ ( posedge clock)
		  ni1i00O62 <= ni1i00O61;
	initial
		ni1i01i67 = 0;
	always @ ( posedge clock)
		  ni1i01i67 <= ni1i01i68;
	event ni1i01i67_event;
	initial
		#1 ->ni1i01i67_event;
	always @(ni1i01i67_event)
		ni1i01i67 <= {1{1'b1}};
	initial
		ni1i01i68 = 0;
	always @ ( posedge clock)
		  ni1i01i68 <= ni1i01i67;
	initial
		ni1i01O65 = 0;
	always @ ( posedge clock)
		  ni1i01O65 <= ni1i01O66;
	event ni1i01O65_event;
	initial
		#1 ->ni1i01O65_event;
	always @(ni1i01O65_event)
		ni1i01O65 <= {1{1'b1}};
	initial
		ni1i01O66 = 0;
	always @ ( posedge clock)
		  ni1i01O66 <= ni1i01O65;
	initial
		ni1i0il59 = 0;
	always @ ( posedge clock)
		  ni1i0il59 <= ni1i0il60;
	event ni1i0il59_event;
	initial
		#1 ->ni1i0il59_event;
	always @(ni1i0il59_event)
		ni1i0il59 <= {1{1'b1}};
	initial
		ni1i0il60 = 0;
	always @ ( posedge clock)
		  ni1i0il60 <= ni1i0il59;
	initial
		ni1i0iO57 = 0;
	always @ ( posedge clock)
		  ni1i0iO57 <= ni1i0iO58;
	event ni1i0iO57_event;
	initial
		#1 ->ni1i0iO57_event;
	always @(ni1i0iO57_event)
		ni1i0iO57 <= {1{1'b1}};
	initial
		ni1i0iO58 = 0;
	always @ ( posedge clock)
		  ni1i0iO58 <= ni1i0iO57;
	initial
		ni1i0ll55 = 0;
	always @ ( posedge clock)
		  ni1i0ll55 <= ni1i0ll56;
	event ni1i0ll55_event;
	initial
		#1 ->ni1i0ll55_event;
	always @(ni1i0ll55_event)
		ni1i0ll55 <= {1{1'b1}};
	initial
		ni1i0ll56 = 0;
	always @ ( posedge clock)
		  ni1i0ll56 <= ni1i0ll55;
	initial
		ni1i0Oi53 = 0;
	always @ ( posedge clock)
		  ni1i0Oi53 <= ni1i0Oi54;
	event ni1i0Oi53_event;
	initial
		#1 ->ni1i0Oi53_event;
	always @(ni1i0Oi53_event)
		ni1i0Oi53 <= {1{1'b1}};
	initial
		ni1i0Oi54 = 0;
	always @ ( posedge clock)
		  ni1i0Oi54 <= ni1i0Oi53;
	initial
		ni1i0Ol51 = 0;
	always @ ( posedge clock)
		  ni1i0Ol51 <= ni1i0Ol52;
	event ni1i0Ol51_event;
	initial
		#1 ->ni1i0Ol51_event;
	always @(ni1i0Ol51_event)
		ni1i0Ol51 <= {1{1'b1}};
	initial
		ni1i0Ol52 = 0;
	always @ ( posedge clock)
		  ni1i0Ol52 <= ni1i0Ol51;
	initial
		ni1i10O79 = 0;
	always @ ( posedge clock)
		  ni1i10O79 <= ni1i10O80;
	event ni1i10O79_event;
	initial
		#1 ->ni1i10O79_event;
	always @(ni1i10O79_event)
		ni1i10O79 <= {1{1'b1}};
	initial
		ni1i10O80 = 0;
	always @ ( posedge clock)
		  ni1i10O80 <= ni1i10O79;
	initial
		ni1i1ii77 = 0;
	always @ ( posedge clock)
		  ni1i1ii77 <= ni1i1ii78;
	event ni1i1ii77_event;
	initial
		#1 ->ni1i1ii77_event;
	always @(ni1i1ii77_event)
		ni1i1ii77 <= {1{1'b1}};
	initial
		ni1i1ii78 = 0;
	always @ ( posedge clock)
		  ni1i1ii78 <= ni1i1ii77;
	initial
		ni1i1li75 = 0;
	always @ ( posedge clock)
		  ni1i1li75 <= ni1i1li76;
	event ni1i1li75_event;
	initial
		#1 ->ni1i1li75_event;
	always @(ni1i1li75_event)
		ni1i1li75 <= {1{1'b1}};
	initial
		ni1i1li76 = 0;
	always @ ( posedge clock)
		  ni1i1li76 <= ni1i1li75;
	initial
		ni1i1ll73 = 0;
	always @ ( posedge clock)
		  ni1i1ll73 <= ni1i1ll74;
	event ni1i1ll73_event;
	initial
		#1 ->ni1i1ll73_event;
	always @(ni1i1ll73_event)
		ni1i1ll73 <= {1{1'b1}};
	initial
		ni1i1ll74 = 0;
	always @ ( posedge clock)
		  ni1i1ll74 <= ni1i1ll73;
	initial
		ni1i1Oi71 = 0;
	always @ ( posedge clock)
		  ni1i1Oi71 <= ni1i1Oi72;
	event ni1i1Oi71_event;
	initial
		#1 ->ni1i1Oi71_event;
	always @(ni1i1Oi71_event)
		ni1i1Oi71 <= {1{1'b1}};
	initial
		ni1i1Oi72 = 0;
	always @ ( posedge clock)
		  ni1i1Oi72 <= ni1i1Oi71;
	initial
		ni1i1Ol69 = 0;
	always @ ( posedge clock)
		  ni1i1Ol69 <= ni1i1Ol70;
	event ni1i1Ol69_event;
	initial
		#1 ->ni1i1Ol69_event;
	always @(ni1i1Ol69_event)
		ni1i1Ol69 <= {1{1'b1}};
	initial
		ni1i1Ol70 = 0;
	always @ ( posedge clock)
		  ni1i1Ol70 <= ni1i1Ol69;
	initial
		ni1ii1i49 = 0;
	always @ ( posedge clock)
		  ni1ii1i49 <= ni1ii1i50;
	event ni1ii1i49_event;
	initial
		#1 ->ni1ii1i49_event;
	always @(ni1ii1i49_event)
		ni1ii1i49 <= {1{1'b1}};
	initial
		ni1ii1i50 = 0;
	always @ ( posedge clock)
		  ni1ii1i50 <= ni1ii1i49;
	initial
		ni1ii1O47 = 0;
	always @ ( posedge clock)
		  ni1ii1O47 <= ni1ii1O48;
	event ni1ii1O47_event;
	initial
		#1 ->ni1ii1O47_event;
	always @(ni1ii1O47_event)
		ni1ii1O47 <= {1{1'b1}};
	initial
		ni1ii1O48 = 0;
	always @ ( posedge clock)
		  ni1ii1O48 <= ni1ii1O47;
	initial
		ni1iill45 = 0;
	always @ ( posedge clock)
		  ni1iill45 <= ni1iill46;
	event ni1iill45_event;
	initial
		#1 ->ni1iill45_event;
	always @(ni1iill45_event)
		ni1iill45 <= {1{1'b1}};
	initial
		ni1iill46 = 0;
	always @ ( posedge clock)
		  ni1iill46 <= ni1iill45;
	initial
		ni1il0i41 = 0;
	always @ ( posedge clock)
		  ni1il0i41 <= ni1il0i42;
	event ni1il0i41_event;
	initial
		#1 ->ni1il0i41_event;
	always @(ni1il0i41_event)
		ni1il0i41 <= {1{1'b1}};
	initial
		ni1il0i42 = 0;
	always @ ( posedge clock)
		  ni1il0i42 <= ni1il0i41;
	initial
		ni1il0l39 = 0;
	always @ ( posedge clock)
		  ni1il0l39 <= ni1il0l40;
	event ni1il0l39_event;
	initial
		#1 ->ni1il0l39_event;
	always @(ni1il0l39_event)
		ni1il0l39 <= {1{1'b1}};
	initial
		ni1il0l40 = 0;
	always @ ( posedge clock)
		  ni1il0l40 <= ni1il0l39;
	initial
		ni1il0O37 = 0;
	always @ ( posedge clock)
		  ni1il0O37 <= ni1il0O38;
	event ni1il0O37_event;
	initial
		#1 ->ni1il0O37_event;
	always @(ni1il0O37_event)
		ni1il0O37 <= {1{1'b1}};
	initial
		ni1il0O38 = 0;
	always @ ( posedge clock)
		  ni1il0O38 <= ni1il0O37;
	initial
		ni1il1O43 = 0;
	always @ ( posedge clock)
		  ni1il1O43 <= ni1il1O44;
	event ni1il1O43_event;
	initial
		#1 ->ni1il1O43_event;
	always @(ni1il1O43_event)
		ni1il1O43 <= {1{1'b1}};
	initial
		ni1il1O44 = 0;
	always @ ( posedge clock)
		  ni1il1O44 <= ni1il1O43;
	initial
		ni1ilii35 = 0;
	always @ ( posedge clock)
		  ni1ilii35 <= ni1ilii36;
	event ni1ilii35_event;
	initial
		#1 ->ni1ilii35_event;
	always @(ni1ilii35_event)
		ni1ilii35 <= {1{1'b1}};
	initial
		ni1ilii36 = 0;
	always @ ( posedge clock)
		  ni1ilii36 <= ni1ilii35;
	initial
		ni1ilil33 = 0;
	always @ ( posedge clock)
		  ni1ilil33 <= ni1ilil34;
	event ni1ilil33_event;
	initial
		#1 ->ni1ilil33_event;
	always @(ni1ilil33_event)
		ni1ilil33 <= {1{1'b1}};
	initial
		ni1ilil34 = 0;
	always @ ( posedge clock)
		  ni1ilil34 <= ni1ilil33;
	initial
		ni1iliO31 = 0;
	always @ ( posedge clock)
		  ni1iliO31 <= ni1iliO32;
	event ni1iliO31_event;
	initial
		#1 ->ni1iliO31_event;
	always @(ni1iliO31_event)
		ni1iliO31 <= {1{1'b1}};
	initial
		ni1iliO32 = 0;
	always @ ( posedge clock)
		  ni1iliO32 <= ni1iliO31;
	initial
		ni1illi29 = 0;
	always @ ( posedge clock)
		  ni1illi29 <= ni1illi30;
	event ni1illi29_event;
	initial
		#1 ->ni1illi29_event;
	always @(ni1illi29_event)
		ni1illi29 <= {1{1'b1}};
	initial
		ni1illi30 = 0;
	always @ ( posedge clock)
		  ni1illi30 <= ni1illi29;
	initial
		ni1illl27 = 0;
	always @ ( posedge clock)
		  ni1illl27 <= ni1illl28;
	event ni1illl27_event;
	initial
		#1 ->ni1illl27_event;
	always @(ni1illl27_event)
		ni1illl27 <= {1{1'b1}};
	initial
		ni1illl28 = 0;
	always @ ( posedge clock)
		  ni1illl28 <= ni1illl27;
	initial
		ni1illO25 = 0;
	always @ ( posedge clock)
		  ni1illO25 <= ni1illO26;
	event ni1illO25_event;
	initial
		#1 ->ni1illO25_event;
	always @(ni1illO25_event)
		ni1illO25 <= {1{1'b1}};
	initial
		ni1illO26 = 0;
	always @ ( posedge clock)
		  ni1illO26 <= ni1illO25;
	initial
		ni1ilOi23 = 0;
	always @ ( posedge clock)
		  ni1ilOi23 <= ni1ilOi24;
	event ni1ilOi23_event;
	initial
		#1 ->ni1ilOi23_event;
	always @(ni1ilOi23_event)
		ni1ilOi23 <= {1{1'b1}};
	initial
		ni1ilOi24 = 0;
	always @ ( posedge clock)
		  ni1ilOi24 <= ni1ilOi23;
	initial
		ni1ilOl21 = 0;
	always @ ( posedge clock)
		  ni1ilOl21 <= ni1ilOl22;
	event ni1ilOl21_event;
	initial
		#1 ->ni1ilOl21_event;
	always @(ni1ilOl21_event)
		ni1ilOl21 <= {1{1'b1}};
	initial
		ni1ilOl22 = 0;
	always @ ( posedge clock)
		  ni1ilOl22 <= ni1ilOl21;
	initial
		ni1ilOO19 = 0;
	always @ ( posedge clock)
		  ni1ilOO19 <= ni1ilOO20;
	event ni1ilOO19_event;
	initial
		#1 ->ni1ilOO19_event;
	always @(ni1ilOO19_event)
		ni1ilOO19 <= {1{1'b1}};
	initial
		ni1ilOO20 = 0;
	always @ ( posedge clock)
		  ni1ilOO20 <= ni1ilOO19;
	initial
		ni1iO0i11 = 0;
	always @ ( posedge clock)
		  ni1iO0i11 <= ni1iO0i12;
	event ni1iO0i11_event;
	initial
		#1 ->ni1iO0i11_event;
	always @(ni1iO0i11_event)
		ni1iO0i11 <= {1{1'b1}};
	initial
		ni1iO0i12 = 0;
	always @ ( posedge clock)
		  ni1iO0i12 <= ni1iO0i11;
	initial
		ni1iO0l10 = 0;
	always @ ( posedge clock)
		  ni1iO0l10 <= ni1iO0l9;
	initial
		ni1iO0l9 = 0;
	always @ ( posedge clock)
		  ni1iO0l9 <= ni1iO0l10;
	event ni1iO0l9_event;
	initial
		#1 ->ni1iO0l9_event;
	always @(ni1iO0l9_event)
		ni1iO0l9 <= {1{1'b1}};
	initial
		ni1iO0O7 = 0;
	always @ ( posedge clock)
		  ni1iO0O7 <= ni1iO0O8;
	event ni1iO0O7_event;
	initial
		#1 ->ni1iO0O7_event;
	always @(ni1iO0O7_event)
		ni1iO0O7 <= {1{1'b1}};
	initial
		ni1iO0O8 = 0;
	always @ ( posedge clock)
		  ni1iO0O8 <= ni1iO0O7;
	initial
		ni1iO1i17 = 0;
	always @ ( posedge clock)
		  ni1iO1i17 <= ni1iO1i18;
	event ni1iO1i17_event;
	initial
		#1 ->ni1iO1i17_event;
	always @(ni1iO1i17_event)
		ni1iO1i17 <= {1{1'b1}};
	initial
		ni1iO1i18 = 0;
	always @ ( posedge clock)
		  ni1iO1i18 <= ni1iO1i17;
	initial
		ni1iO1l15 = 0;
	always @ ( posedge clock)
		  ni1iO1l15 <= ni1iO1l16;
	event ni1iO1l15_event;
	initial
		#1 ->ni1iO1l15_event;
	always @(ni1iO1l15_event)
		ni1iO1l15 <= {1{1'b1}};
	initial
		ni1iO1l16 = 0;
	always @ ( posedge clock)
		  ni1iO1l16 <= ni1iO1l15;
	initial
		ni1iO1O13 = 0;
	always @ ( posedge clock)
		  ni1iO1O13 <= ni1iO1O14;
	event ni1iO1O13_event;
	initial
		#1 ->ni1iO1O13_event;
	always @(ni1iO1O13_event)
		ni1iO1O13 <= {1{1'b1}};
	initial
		ni1iO1O14 = 0;
	always @ ( posedge clock)
		  ni1iO1O14 <= ni1iO1O13;
	initial
		ni1iOii5 = 0;
	always @ ( posedge clock)
		  ni1iOii5 <= ni1iOii6;
	event ni1iOii5_event;
	initial
		#1 ->ni1iOii5_event;
	always @(ni1iOii5_event)
		ni1iOii5 <= {1{1'b1}};
	initial
		ni1iOii6 = 0;
	always @ ( posedge clock)
		  ni1iOii6 <= ni1iOii5;
	initial
		ni1iOil3 = 0;
	always @ ( posedge clock)
		  ni1iOil3 <= ni1iOil4;
	event ni1iOil3_event;
	initial
		#1 ->ni1iOil3_event;
	always @(ni1iOil3_event)
		ni1iOil3 <= {1{1'b1}};
	initial
		ni1iOil4 = 0;
	always @ ( posedge clock)
		  ni1iOil4 <= ni1iOil3;
	initial
		ni1iOll1 = 0;
	always @ ( posedge clock)
		  ni1iOll1 <= ni1iOll2;
	event ni1iOll1_event;
	initial
		#1 ->ni1iOll1_event;
	always @(ni1iOll1_event)
		ni1iOll1 <= {1{1'b1}};
	initial
		ni1iOll2 = 0;
	always @ ( posedge clock)
		  ni1iOll2 <= ni1iOll1;
	initial
	begin
		n100i = 0;
		n100l = 0;
		n100O = 0;
		n101i = 0;
		n101l = 0;
		n101O = 0;
		n10ii = 0;
		n10il = 0;
		n10iO = 0;
		n10li = 0;
		n10ll = 0;
		n10lO = 0;
		n10Oi = 0;
		n10Ol = 0;
		n10OO = 0;
		n110i = 0;
		n110l = 0;
		n110O = 0;
		n111i = 0;
		n111l = 0;
		n111O = 0;
		n11ii = 0;
		n11il = 0;
		n11iO = 0;
		n11li = 0;
		n11ll = 0;
		n11lO = 0;
		n11Oi = 0;
		n11Ol = 0;
		n11OO = 0;
		n1i0i = 0;
		n1i0l = 0;
		n1i0O = 0;
		n1i1i = 0;
		n1i1l = 0;
		n1i1O = 0;
		n1iii = 0;
		n1iil = 0;
		n1ili = 0;
		nlO10l = 0;
		nlOOOi = 0;
		nlOOOl = 0;
		nlOOOO = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			n100i <= 0;
			n100l <= 0;
			n100O <= 0;
			n101i <= 0;
			n101l <= 0;
			n101O <= 0;
			n10ii <= 0;
			n10il <= 0;
			n10iO <= 0;
			n10li <= 0;
			n10ll <= 0;
			n10lO <= 0;
			n10Oi <= 0;
			n10Ol <= 0;
			n10OO <= 0;
			n110i <= 0;
			n110l <= 0;
			n110O <= 0;
			n111i <= 0;
			n111l <= 0;
			n111O <= 0;
			n11ii <= 0;
			n11il <= 0;
			n11iO <= 0;
			n11li <= 0;
			n11ll <= 0;
			n11lO <= 0;
			n11Oi <= 0;
			n11Ol <= 0;
			n11OO <= 0;
			n1i0i <= 0;
			n1i0l <= 0;
			n1i0O <= 0;
			n1i1i <= 0;
			n1i1l <= 0;
			n1i1O <= 0;
			n1iii <= 0;
			n1iil <= 0;
			n1ili <= 0;
			nlO10l <= 0;
			nlOOOi <= 0;
			nlOOOl <= 0;
			nlOOOO <= 0;
		end
		else if  (ni1iiOO == 1'b1) 
		begin
			n100i <= wire_n1O0i_o;
			n100l <= wire_n1O0l_o;
			n100O <= wire_n1O0O_o;
			n101i <= wire_n1O1i_o;
			n101l <= wire_n1O1l_o;
			n101O <= wire_n1O1O_o;
			n10ii <= wire_n1Oii_o;
			n10il <= wire_n1Oil_o;
			n10iO <= wire_n1OiO_o;
			n10li <= wire_n1Oli_o;
			n10ll <= wire_n1Oll_o;
			n10lO <= wire_n1OlO_o;
			n10Oi <= wire_n1OOi_o;
			n10Ol <= wire_n1OOl_o;
			n10OO <= wire_n1OOO_o;
			n110i <= wire_n1l0i_o;
			n110l <= wire_n1l0l_o;
			n110O <= wire_n1l0O_o;
			n111i <= wire_n1l1i_o;
			n111l <= wire_n1l1l_o;
			n111O <= wire_n1l1O_o;
			n11ii <= wire_n1lii_o;
			n11il <= wire_n1lil_o;
			n11iO <= wire_n1liO_o;
			n11li <= wire_n1lli_o;
			n11ll <= wire_n1lll_o;
			n11lO <= wire_n1llO_o;
			n11Oi <= wire_n1lOi_o;
			n11Ol <= wire_n1lOl_o;
			n11OO <= wire_n1lOO_o;
			n1i0i <= wire_nl001iO_q[1];
			n1i0l <= wire_nl001iO_q[2];
			n1i0O <= wire_nl001iO_q[3];
			n1i1i <= wire_n011i_o;
			n1i1l <= wire_n011l_o;
			n1i1O <= wire_nl001iO_q[0];
			n1iii <= wire_nl001iO_q[4];
			n1iil <= wire_nl001iO_q[5];
			n1ili <= wire_nl001iO_q[6];
			nlO10l <= wire_n1ilO_o;
			nlOOOi <= wire_n1iOi_o;
			nlOOOl <= wire_n1iOl_o;
			nlOOOO <= wire_n1iOO_o;
		end
	end
	initial
	begin
		ni0101l = 0;
		ni01lil = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			ni0101l <= 0;
			ni01lil <= 0;
		end
		else if  (n0OOOil == 1'b0) 
		begin
			ni0101l <= n0OOOii;
			ni01lil <= n0OOOii;
		end
	end
	initial
	begin
		n000i = 0;
		n000l = 0;
		n000O = 0;
		n001i = 0;
		n001l = 0;
		n001O = 0;
		n00ii = 0;
		n00il = 0;
		n00iO = 0;
		n00li = 0;
		n00ll = 0;
		n00lO = 0;
		n00Oi = 0;
		n00Ol = 0;
		n00OO = 0;
		n010i = 0;
		n010l = 0;
		n010O = 0;
		n011O = 0;
		n01ii = 0;
		n01il = 0;
		n01iO = 0;
		n01li = 0;
		n01ll = 0;
		n01lO = 0;
		n01Oi = 0;
		n01Ol = 0;
		n01OO = 0;
		n0i0i = 0;
		n0i0l = 0;
		n0i0O = 0;
		n0i1i = 0;
		n0i1l = 0;
		n0i1O = 0;
		n0iii = 0;
		n0iil = 0;
		n0iiO = 0;
		n0ili = 0;
		n0ill = 0;
		n0ilO = 0;
		n0iOi = 0;
		n0iOl = 0;
		n0iOO = 0;
		n0l0i = 0;
		n0l0l = 0;
		n0l0O = 0;
		n0l1i = 0;
		n0l1l = 0;
		n0l1O = 0;
		n0lii = 0;
		n0lil = 0;
		n0liO = 0;
		n0lli = 0;
		n0lll = 0;
		n0llO = 0;
		n0lOi = 0;
		n0lOl = 0;
		n0lOO = 0;
		n0O0i = 0;
		n0O0l = 0;
		n0O0O = 0;
		n0O1i = 0;
		n0O1l = 0;
		n0O1O = 0;
		n0Oii = 0;
		n0Oil = 0;
		n0OiO = 0;
		n0Oli = 0;
		n0Oll = 0;
		n0OlO = 0;
		n0OOi = 0;
		n0OOl = 0;
		n0OOO = 0;
		n1ill = 0;
		ni10l = 0;
		ni11i = 0;
		ni11l = 0;
		ni11O = 0;
	end
	always @ (clock or wire_ni10i_PRN or wire_ni10i_CLRN)
	begin
		if (wire_ni10i_PRN == 1'b0) 
		begin
			n000i <= 1;
			n000l <= 1;
			n000O <= 1;
			n001i <= 1;
			n001l <= 1;
			n001O <= 1;
			n00ii <= 1;
			n00il <= 1;
			n00iO <= 1;
			n00li <= 1;
			n00ll <= 1;
			n00lO <= 1;
			n00Oi <= 1;
			n00Ol <= 1;
			n00OO <= 1;
			n010i <= 1;
			n010l <= 1;
			n010O <= 1;
			n011O <= 1;
			n01ii <= 1;
			n01il <= 1;
			n01iO <= 1;
			n01li <= 1;
			n01ll <= 1;
			n01lO <= 1;
			n01Oi <= 1;
			n01Ol <= 1;
			n01OO <= 1;
			n0i0i <= 1;
			n0i0l <= 1;
			n0i0O <= 1;
			n0i1i <= 1;
			n0i1l <= 1;
			n0i1O <= 1;
			n0iii <= 1;
			n0iil <= 1;
			n0iiO <= 1;
			n0ili <= 1;
			n0ill <= 1;
			n0ilO <= 1;
			n0iOi <= 1;
			n0iOl <= 1;
			n0iOO <= 1;
			n0l0i <= 1;
			n0l0l <= 1;
			n0l0O <= 1;
			n0l1i <= 1;
			n0l1l <= 1;
			n0l1O <= 1;
			n0lii <= 1;
			n0lil <= 1;
			n0liO <= 1;
			n0lli <= 1;
			n0lll <= 1;
			n0llO <= 1;
			n0lOi <= 1;
			n0lOl <= 1;
			n0lOO <= 1;
			n0O0i <= 1;
			n0O0l <= 1;
			n0O0O <= 1;
			n0O1i <= 1;
			n0O1l <= 1;
			n0O1O <= 1;
			n0Oii <= 1;
			n0Oil <= 1;
			n0OiO <= 1;
			n0Oli <= 1;
			n0Oll <= 1;
			n0OlO <= 1;
			n0OOi <= 1;
			n0OOl <= 1;
			n0OOO <= 1;
			n1ill <= 1;
			ni10l <= 1;
			ni11i <= 1;
			ni11l <= 1;
			ni11O <= 1;
		end
		else if  (wire_ni10i_CLRN == 1'b0) 
		begin
			n000i <= 0;
			n000l <= 0;
			n000O <= 0;
			n001i <= 0;
			n001l <= 0;
			n001O <= 0;
			n00ii <= 0;
			n00il <= 0;
			n00iO <= 0;
			n00li <= 0;
			n00ll <= 0;
			n00lO <= 0;
			n00Oi <= 0;
			n00Ol <= 0;
			n00OO <= 0;
			n010i <= 0;
			n010l <= 0;
			n010O <= 0;
			n011O <= 0;
			n01ii <= 0;
			n01il <= 0;
			n01iO <= 0;
			n01li <= 0;
			n01ll <= 0;
			n01lO <= 0;
			n01Oi <= 0;
			n01Ol <= 0;
			n01OO <= 0;
			n0i0i <= 0;
			n0i0l <= 0;
			n0i0O <= 0;
			n0i1i <= 0;
			n0i1l <= 0;
			n0i1O <= 0;
			n0iii <= 0;
			n0iil <= 0;
			n0iiO <= 0;
			n0ili <= 0;
			n0ill <= 0;
			n0ilO <= 0;
			n0iOi <= 0;
			n0iOl <= 0;
			n0iOO <= 0;
			n0l0i <= 0;
			n0l0l <= 0;
			n0l0O <= 0;
			n0l1i <= 0;
			n0l1l <= 0;
			n0l1O <= 0;
			n0lii <= 0;
			n0lil <= 0;
			n0liO <= 0;
			n0lli <= 0;
			n0lll <= 0;
			n0llO <= 0;
			n0lOi <= 0;
			n0lOl <= 0;
			n0lOO <= 0;
			n0O0i <= 0;
			n0O0l <= 0;
			n0O0O <= 0;
			n0O1i <= 0;
			n0O1l <= 0;
			n0O1O <= 0;
			n0Oii <= 0;
			n0Oil <= 0;
			n0OiO <= 0;
			n0Oli <= 0;
			n0Oll <= 0;
			n0OlO <= 0;
			n0OOi <= 0;
			n0OOl <= 0;
			n0OOO <= 0;
			n1ill <= 0;
			ni10l <= 0;
			ni11i <= 0;
			ni11l <= 0;
			ni11O <= 0;
		end
		else if  (ni1il1l == 1'b1) 
		if (clock != ni10i_clk_prev && clock == 1'b1) 
		begin
			n000i <= wire_ni0il_o;
			n000l <= wire_ni0iO_o;
			n000O <= wire_ni0li_o;
			n001i <= wire_ni00l_o;
			n001l <= wire_ni00O_o;
			n001O <= wire_ni0ii_o;
			n00ii <= wire_ni0ll_o;
			n00il <= wire_ni0lO_o;
			n00iO <= wire_ni0Oi_o;
			n00li <= wire_ni0Ol_o;
			n00ll <= wire_ni0OO_o;
			n00lO <= wire_nii1i_o;
			n00Oi <= wire_nii1l_o;
			n00Ol <= wire_nii1O_o;
			n00OO <= wire_nii0i_o;
			n010i <= wire_ni1il_o;
			n010l <= wire_ni1iO_o;
			n010O <= wire_ni1li_o;
			n011O <= wire_ni1ii_o;
			n01ii <= wire_ni1ll_o;
			n01il <= wire_ni1lO_o;
			n01iO <= wire_ni1Oi_o;
			n01li <= wire_ni1Ol_o;
			n01ll <= wire_ni1OO_o;
			n01lO <= wire_ni01i_o;
			n01Oi <= wire_ni01l_o;
			n01Ol <= wire_ni01O_o;
			n01OO <= wire_ni00i_o;
			n0i0i <= wire_niiil_o;
			n0i0l <= wire_niiiO_o;
			n0i0O <= wire_niili_o;
			n0i1i <= wire_nii0l_o;
			n0i1l <= wire_nii0O_o;
			n0i1O <= wire_niiii_o;
			n0iii <= wire_niill_o;
			n0iil <= wire_niilO_o;
			n0iiO <= wire_niiOi_o;
			n0ili <= wire_niiOl_o;
			n0ill <= wire_niiOO_o;
			n0ilO <= wire_nil1i_o;
			n0iOi <= wire_nil1l_o;
			n0iOl <= wire_nil1O_o;
			n0iOO <= wire_nil0i_o;
			n0l0i <= wire_nilil_o;
			n0l0l <= wire_niliO_o;
			n0l0O <= wire_nilli_o;
			n0l1i <= wire_nil0l_o;
			n0l1l <= wire_nil0O_o;
			n0l1O <= wire_nilii_o;
			n0lii <= wire_nilll_o;
			n0lil <= wire_nillO_o;
			n0liO <= wire_nilOi_o;
			n0lli <= wire_nilOl_o;
			n0lll <= wire_nilOO_o;
			n0llO <= wire_niO1i_o;
			n0lOi <= wire_niO1l_o;
			n0lOl <= wire_niO1O_o;
			n0lOO <= wire_niO0i_o;
			n0O0i <= wire_niOil_o;
			n0O0l <= wire_niOiO_o;
			n0O0O <= ni11O;
			n0O1i <= wire_niO0l_o;
			n0O1l <= wire_niO0O_o;
			n0O1O <= wire_niOii_o;
			n0Oii <= wire_niOli_o;
			n0Oil <= wire_niOll_o;
			n0OiO <= wire_niOlO_o;
			n0Oli <= wire_niOOi_o;
			n0Oll <= wire_niOOl_o;
			n0OlO <= wire_nl01O0i_q[0];
			n0OOi <= wire_nl01O0i_q[1];
			n0OOl <= wire_nl01O0i_q[2];
			n0OOO <= wire_nl01O0i_q[3];
			n1ill <= wire_ni10O_o;
			ni10l <= wire_nl01O0i_q[7];
			ni11i <= wire_nl01O0i_q[4];
			ni11l <= wire_nl01O0i_q[5];
			ni11O <= wire_nl01O0i_q[6];
		end
		ni10i_clk_prev <= clock;
	end
	assign
		wire_ni10i_CLRN = ((ni1il0i42 ^ ni1il0i41) & (~ reset)),
		wire_ni10i_PRN = (ni1il1O44 ^ ni1il1O43);
	event n000i_event;
	event n000l_event;
	event n000O_event;
	event n001i_event;
	event n001l_event;
	event n001O_event;
	event n00ii_event;
	event n00il_event;
	event n00iO_event;
	event n00li_event;
	event n00ll_event;
	event n00lO_event;
	event n00Oi_event;
	event n00Ol_event;
	event n00OO_event;
	event n010i_event;
	event n010l_event;
	event n010O_event;
	event n011O_event;
	event n01ii_event;
	event n01il_event;
	event n01iO_event;
	event n01li_event;
	event n01ll_event;
	event n01lO_event;
	event n01Oi_event;
	event n01Ol_event;
	event n01OO_event;
	event n0i0i_event;
	event n0i0l_event;
	event n0i0O_event;
	event n0i1i_event;
	event n0i1l_event;
	event n0i1O_event;
	event n0iii_event;
	event n0iil_event;
	event n0iiO_event;
	event n0ili_event;
	event n0ill_event;
	event n0ilO_event;
	event n0iOi_event;
	event n0iOl_event;
	event n0iOO_event;
	event n0l0i_event;
	event n0l0l_event;
	event n0l0O_event;
	event n0l1i_event;
	event n0l1l_event;
	event n0l1O_event;
	event n0lii_event;
	event n0lil_event;
	event n0liO_event;
	event n0lli_event;
	event n0lll_event;
	event n0llO_event;
	event n0lOi_event;
	event n0lOl_event;
	event n0lOO_event;
	event n0O0i_event;
	event n0O0l_event;
	event n0O0O_event;
	event n0O1i_event;
	event n0O1l_event;
	event n0O1O_event;
	event n0Oii_event;
	event n0Oil_event;
	event n0OiO_event;
	event n0Oli_event;
	event n0Oll_event;
	event n0OlO_event;
	event n0OOi_event;
	event n0OOl_event;
	event n0OOO_event;
	event n1ill_event;
	event ni10l_event;
	event ni11i_event;
	event ni11l_event;
	event ni11O_event;
	initial
		#1 ->n000i_event;
	initial
		#1 ->n000l_event;
	initial
		#1 ->n000O_event;
	initial
		#1 ->n001i_event;
	initial
		#1 ->n001l_event;
	initial
		#1 ->n001O_event;
	initial
		#1 ->n00ii_event;
	initial
		#1 ->n00il_event;
	initial
		#1 ->n00iO_event;
	initial
		#1 ->n00li_event;
	initial
		#1 ->n00ll_event;
	initial
		#1 ->n00lO_event;
	initial
		#1 ->n00Oi_event;
	initial
		#1 ->n00Ol_event;
	initial
		#1 ->n00OO_event;
	initial
		#1 ->n010i_event;
	initial
		#1 ->n010l_event;
	initial
		#1 ->n010O_event;
	initial
		#1 ->n011O_event;
	initial
		#1 ->n01ii_event;
	initial
		#1 ->n01il_event;
	initial
		#1 ->n01iO_event;
	initial
		#1 ->n01li_event;
	initial
		#1 ->n01ll_event;
	initial
		#1 ->n01lO_event;
	initial
		#1 ->n01Oi_event;
	initial
		#1 ->n01Ol_event;
	initial
		#1 ->n01OO_event;
	initial
		#1 ->n0i0i_event;
	initial
		#1 ->n0i0l_event;
	initial
		#1 ->n0i0O_event;
	initial
		#1 ->n0i1i_event;
	initial
		#1 ->n0i1l_event;
	initial
		#1 ->n0i1O_event;
	initial
		#1 ->n0iii_event;
	initial
		#1 ->n0iil_event;
	initial
		#1 ->n0iiO_event;
	initial
		#1 ->n0ili_event;
	initial
		#1 ->n0ill_event;
	initial
		#1 ->n0ilO_event;
	initial
		#1 ->n0iOi_event;
	initial
		#1 ->n0iOl_event;
	initial
		#1 ->n0iOO_event;
	initial
		#1 ->n0l0i_event;
	initial
		#1 ->n0l0l_event;
	initial
		#1 ->n0l0O_event;
	initial
		#1 ->n0l1i_event;
	initial
		#1 ->n0l1l_event;
	initial
		#1 ->n0l1O_event;
	initial
		#1 ->n0lii_event;
	initial
		#1 ->n0lil_event;
	initial
		#1 ->n0liO_event;
	initial
		#1 ->n0lli_event;
	initial
		#1 ->n0lll_event;
	initial
		#1 ->n0llO_event;
	initial
		#1 ->n0lOi_event;
	initial
		#1 ->n0lOl_event;
	initial
		#1 ->n0lOO_event;
	initial
		#1 ->n0O0i_event;
	initial
		#1 ->n0O0l_event;
	initial
		#1 ->n0O0O_event;
	initial
		#1 ->n0O1i_event;
	initial
		#1 ->n0O1l_event;
	initial
		#1 ->n0O1O_event;
	initial
		#1 ->n0Oii_event;
	initial
		#1 ->n0Oil_event;
	initial
		#1 ->n0OiO_event;
	initial
		#1 ->n0Oli_event;
	initial
		#1 ->n0Oll_event;
	initial
		#1 ->n0OlO_event;
	initial
		#1 ->n0OOi_event;
	initial
		#1 ->n0OOl_event;
	initial
		#1 ->n0OOO_event;
	initial
		#1 ->n1ill_event;
	initial
		#1 ->ni10l_event;
	initial
		#1 ->ni11i_event;
	initial
		#1 ->ni11l_event;
	initial
		#1 ->ni11O_event;
	always @(n000i_event)
		n000i <= 1;
	always @(n000l_event)
		n000l <= 1;
	always @(n000O_event)
		n000O <= 1;
	always @(n001i_event)
		n001i <= 1;
	always @(n001l_event)
		n001l <= 1;
	always @(n001O_event)
		n001O <= 1;
	always @(n00ii_event)
		n00ii <= 1;
	always @(n00il_event)
		n00il <= 1;
	always @(n00iO_event)
		n00iO <= 1;
	always @(n00li_event)
		n00li <= 1;
	always @(n00ll_event)
		n00ll <= 1;
	always @(n00lO_event)
		n00lO <= 1;
	always @(n00Oi_event)
		n00Oi <= 1;
	always @(n00Ol_event)
		n00Ol <= 1;
	always @(n00OO_event)
		n00OO <= 1;
	always @(n010i_event)
		n010i <= 1;
	always @(n010l_event)
		n010l <= 1;
	always @(n010O_event)
		n010O <= 1;
	always @(n011O_event)
		n011O <= 1;
	always @(n01ii_event)
		n01ii <= 1;
	always @(n01il_event)
		n01il <= 1;
	always @(n01iO_event)
		n01iO <= 1;
	always @(n01li_event)
		n01li <= 1;
	always @(n01ll_event)
		n01ll <= 1;
	always @(n01lO_event)
		n01lO <= 1;
	always @(n01Oi_event)
		n01Oi <= 1;
	always @(n01Ol_event)
		n01Ol <= 1;
	always @(n01OO_event)
		n01OO <= 1;
	always @(n0i0i_event)
		n0i0i <= 1;
	always @(n0i0l_event)
		n0i0l <= 1;
	always @(n0i0O_event)
		n0i0O <= 1;
	always @(n0i1i_event)
		n0i1i <= 1;
	always @(n0i1l_event)
		n0i1l <= 1;
	always @(n0i1O_event)
		n0i1O <= 1;
	always @(n0iii_event)
		n0iii <= 1;
	always @(n0iil_event)
		n0iil <= 1;
	always @(n0iiO_event)
		n0iiO <= 1;
	always @(n0ili_event)
		n0ili <= 1;
	always @(n0ill_event)
		n0ill <= 1;
	always @(n0ilO_event)
		n0ilO <= 1;
	always @(n0iOi_event)
		n0iOi <= 1;
	always @(n0iOl_event)
		n0iOl <= 1;
	always @(n0iOO_event)
		n0iOO <= 1;
	always @(n0l0i_event)
		n0l0i <= 1;
	always @(n0l0l_event)
		n0l0l <= 1;
	always @(n0l0O_event)
		n0l0O <= 1;
	always @(n0l1i_event)
		n0l1i <= 1;
	always @(n0l1l_event)
		n0l1l <= 1;
	always @(n0l1O_event)
		n0l1O <= 1;
	always @(n0lii_event)
		n0lii <= 1;
	always @(n0lil_event)
		n0lil <= 1;
	always @(n0liO_event)
		n0liO <= 1;
	always @(n0lli_event)
		n0lli <= 1;
	always @(n0lll_event)
		n0lll <= 1;
	always @(n0llO_event)
		n0llO <= 1;
	always @(n0lOi_event)
		n0lOi <= 1;
	always @(n0lOl_event)
		n0lOl <= 1;
	always @(n0lOO_event)
		n0lOO <= 1;
	always @(n0O0i_event)
		n0O0i <= 1;
	always @(n0O0l_event)
		n0O0l <= 1;
	always @(n0O0O_event)
		n0O0O <= 1;
	always @(n0O1i_event)
		n0O1i <= 1;
	always @(n0O1l_event)
		n0O1l <= 1;
	always @(n0O1O_event)
		n0O1O <= 1;
	always @(n0Oii_event)
		n0Oii <= 1;
	always @(n0Oil_event)
		n0Oil <= 1;
	always @(n0OiO_event)
		n0OiO <= 1;
	always @(n0Oli_event)
		n0Oli <= 1;
	always @(n0Oll_event)
		n0Oll <= 1;
	always @(n0OlO_event)
		n0OlO <= 1;
	always @(n0OOi_event)
		n0OOi <= 1;
	always @(n0OOl_event)
		n0OOl <= 1;
	always @(n0OOO_event)
		n0OOO <= 1;
	always @(n1ill_event)
		n1ill <= 1;
	always @(ni10l_event)
		ni10l <= 1;
	always @(ni11i_event)
		ni11i <= 1;
	always @(ni11l_event)
		ni11l <= 1;
	always @(ni11O_event)
		ni11O <= 1;
	initial
	begin
		nii010i = 0;
		nii010l = 0;
		nii010O = 0;
		nii01ii = 0;
		nii01il = 0;
		nii01li = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nii010i <= 0;
			nii010l <= 0;
			nii010O <= 0;
			nii01ii <= 0;
			nii01il <= 0;
			nii01li <= 0;
		end
		else if  (ni1111O == 1'b1) 
		begin
			nii010i <= wire_nii01lO_dataout;
			nii010l <= wire_nii01Oi_dataout;
			nii010O <= wire_nii01Ol_dataout;
			nii01ii <= wire_nii01OO_dataout;
			nii01il <= wire_nii001i_dataout;
			nii01li <= wire_nii01ll_dataout;
		end
	end
	initial
	begin
		nii00li = 0;
		nii0i0i = 0;
		nii0i0l = 0;
		nii0i0O = 0;
		nii0i1i = 0;
		nii0i1l = 0;
		nii0i1O = 0;
		nii0iii = 0;
		nii0iil = 0;
		nii0iiO = 0;
		nii0ili = 0;
		nii0ill = 0;
		nii0ilO = 0;
		nii0iOi = 0;
		nii0iOl = 0;
		nii0iOO = 0;
		nii0l0i = 0;
		nii0l0l = 0;
		nii0l0O = 0;
		nii0l1i = 0;
		nii0l1l = 0;
		nii0l1O = 0;
		nii0lii = 0;
		nii0lil = 0;
		nii0lli = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nii00li <= 0;
			nii0i0i <= 0;
			nii0i0l <= 0;
			nii0i0O <= 0;
			nii0i1i <= 0;
			nii0i1l <= 0;
			nii0i1O <= 0;
			nii0iii <= 0;
			nii0iil <= 0;
			nii0iiO <= 0;
			nii0ili <= 0;
			nii0ill <= 0;
			nii0ilO <= 0;
			nii0iOi <= 0;
			nii0iOl <= 0;
			nii0iOO <= 0;
			nii0l0i <= 0;
			nii0l0l <= 0;
			nii0l0O <= 0;
			nii0l1i <= 0;
			nii0l1l <= 0;
			nii0l1O <= 0;
			nii0lii <= 0;
			nii0lil <= 0;
			nii0lli <= 0;
		end
		else if  (ni111ii == 1'b1) 
		begin
			nii00li <= wire_niiOl0l_dataout;
			nii0i0i <= wire_niiO0Ol_dataout;
			nii0i0l <= wire_niiO0OO_dataout;
			nii0i0O <= wire_niiOi1i_dataout;
			nii0i1i <= wire_niiO0ll_dataout;
			nii0i1l <= wire_niiO0lO_dataout;
			nii0i1O <= wire_niiO0Oi_dataout;
			nii0iii <= wire_niiOi1l_dataout;
			nii0iil <= wire_niiOi1O_dataout;
			nii0iiO <= wire_niiOi0i_dataout;
			nii0ili <= wire_niiOi0l_dataout;
			nii0ill <= wire_niiOi0O_dataout;
			nii0ilO <= wire_niiOiii_dataout;
			nii0iOi <= wire_niiOiil_dataout;
			nii0iOl <= wire_niiOiiO_dataout;
			nii0iOO <= wire_niiOili_dataout;
			nii0l0i <= wire_niiOiOl_dataout;
			nii0l0l <= wire_niiOiOO_dataout;
			nii0l0O <= wire_niiOl1i_dataout;
			nii0l1i <= wire_niiOill_dataout;
			nii0l1l <= wire_niiOilO_dataout;
			nii0l1O <= wire_niiOiOi_dataout;
			nii0lii <= wire_niiOl1l_dataout;
			nii0lil <= wire_niiOl1O_dataout;
			nii0lli <= wire_niiOl0i_dataout;
		end
	end
	initial
	begin
		ni0O00i = 0;
		ni0O00l = 0;
		ni0O00O = 0;
		ni0O01i = 0;
		ni0O01l = 0;
		ni0O01O = 0;
		ni0O0ii = 0;
		ni0O0il = 0;
		ni0O0iO = 0;
		ni0O0li = 0;
		ni0O0ll = 0;
		ni0O0lO = 0;
		ni0O0Oi = 0;
		ni0O0Ol = 0;
		ni0O0OO = 0;
		ni0O1iO = 0;
		ni0O1li = 0;
		ni0O1ll = 0;
		ni0O1lO = 0;
		ni0O1Oi = 0;
		ni0O1Ol = 0;
		ni0O1OO = 0;
		ni0Oi0l = 0;
		ni0Oi1i = 0;
		ni0Oi1l = 0;
		nii110i = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			ni0O00i <= 0;
			ni0O00l <= 0;
			ni0O00O <= 0;
			ni0O01i <= 0;
			ni0O01l <= 0;
			ni0O01O <= 0;
			ni0O0ii <= 0;
			ni0O0il <= 0;
			ni0O0iO <= 0;
			ni0O0li <= 0;
			ni0O0ll <= 0;
			ni0O0lO <= 0;
			ni0O0Oi <= 0;
			ni0O0Ol <= 0;
			ni0O0OO <= 0;
			ni0O1iO <= 0;
			ni0O1li <= 0;
			ni0O1ll <= 0;
			ni0O1lO <= 0;
			ni0O1Oi <= 0;
			ni0O1Ol <= 0;
			ni0O1OO <= 0;
			ni0Oi0l <= 0;
			ni0Oi1i <= 0;
			ni0Oi1l <= 0;
			nii110i <= 0;
		end
		else if  (ni1iiii == 1'b0) 
		begin
			ni0O00i <= wire_ni0Olil_dataout;
			ni0O00l <= wire_ni0OliO_dataout;
			ni0O00O <= wire_ni0Olli_dataout;
			ni0O01i <= wire_ni0Ol0l_dataout;
			ni0O01l <= wire_ni0Ol0O_dataout;
			ni0O01O <= wire_ni0Olii_dataout;
			ni0O0ii <= wire_ni0Olll_dataout;
			ni0O0il <= wire_ni0OllO_dataout;
			ni0O0iO <= wire_ni0OlOi_dataout;
			ni0O0li <= wire_ni0OlOl_dataout;
			ni0O0ll <= wire_ni0OlOO_dataout;
			ni0O0lO <= wire_ni0OO1i_dataout;
			ni0O0Oi <= wire_ni0OO1l_dataout;
			ni0O0Ol <= wire_ni0OO1O_dataout;
			ni0O0OO <= wire_ni0OO0i_dataout;
			ni0O1iO <= wire_ni0OiOi_dataout;
			ni0O1li <= wire_ni0OiOl_dataout;
			ni0O1ll <= wire_ni0OiOO_dataout;
			ni0O1lO <= wire_ni0Ol1i_dataout;
			ni0O1Oi <= wire_ni0Ol1l_dataout;
			ni0O1Ol <= wire_ni0Ol1O_dataout;
			ni0O1OO <= wire_ni0Ol0i_dataout;
			ni0Oi0l <= wire_ni011Ol_o;
			ni0Oi1i <= wire_ni0OO0l_dataout;
			ni0Oi1l <= wire_ni0OO0O_dataout;
			nii110i <= wire_ni0OilO_dataout;
		end
	end
	event ni0O00i_event;
	event ni0O00l_event;
	event ni0O00O_event;
	event ni0O01i_event;
	event ni0O01l_event;
	event ni0O01O_event;
	event ni0O0ii_event;
	event ni0O0il_event;
	event ni0O0iO_event;
	event ni0O0li_event;
	event ni0O0ll_event;
	event ni0O0lO_event;
	event ni0O0Oi_event;
	event ni0O0Ol_event;
	event ni0O0OO_event;
	event ni0O1iO_event;
	event ni0O1li_event;
	event ni0O1ll_event;
	event ni0O1lO_event;
	event ni0O1Oi_event;
	event ni0O1Ol_event;
	event ni0O1OO_event;
	event ni0Oi0l_event;
	event ni0Oi1i_event;
	event ni0Oi1l_event;
	event nii110i_event;
	initial
		#1 ->ni0O00i_event;
	initial
		#1 ->ni0O00l_event;
	initial
		#1 ->ni0O00O_event;
	initial
		#1 ->ni0O01i_event;
	initial
		#1 ->ni0O01l_event;
	initial
		#1 ->ni0O01O_event;
	initial
		#1 ->ni0O0ii_event;
	initial
		#1 ->ni0O0il_event;
	initial
		#1 ->ni0O0iO_event;
	initial
		#1 ->ni0O0li_event;
	initial
		#1 ->ni0O0ll_event;
	initial
		#1 ->ni0O0lO_event;
	initial
		#1 ->ni0O0Oi_event;
	initial
		#1 ->ni0O0Ol_event;
	initial
		#1 ->ni0O0OO_event;
	initial
		#1 ->ni0O1iO_event;
	initial
		#1 ->ni0O1li_event;
	initial
		#1 ->ni0O1ll_event;
	initial
		#1 ->ni0O1lO_event;
	initial
		#1 ->ni0O1Oi_event;
	initial
		#1 ->ni0O1Ol_event;
	initial
		#1 ->ni0O1OO_event;
	initial
		#1 ->ni0Oi0l_event;
	initial
		#1 ->ni0Oi1i_event;
	initial
		#1 ->ni0Oi1l_event;
	initial
		#1 ->nii110i_event;
	always @(ni0O00i_event)
		ni0O00i <= 1;
	always @(ni0O00l_event)
		ni0O00l <= 1;
	always @(ni0O00O_event)
		ni0O00O <= 1;
	always @(ni0O01i_event)
		ni0O01i <= 1;
	always @(ni0O01l_event)
		ni0O01l <= 1;
	always @(ni0O01O_event)
		ni0O01O <= 1;
	always @(ni0O0ii_event)
		ni0O0ii <= 1;
	always @(ni0O0il_event)
		ni0O0il <= 1;
	always @(ni0O0iO_event)
		ni0O0iO <= 1;
	always @(ni0O0li_event)
		ni0O0li <= 1;
	always @(ni0O0ll_event)
		ni0O0ll <= 1;
	always @(ni0O0lO_event)
		ni0O0lO <= 1;
	always @(ni0O0Oi_event)
		ni0O0Oi <= 1;
	always @(ni0O0Ol_event)
		ni0O0Ol <= 1;
	always @(ni0O0OO_event)
		ni0O0OO <= 1;
	always @(ni0O1iO_event)
		ni0O1iO <= 1;
	always @(ni0O1li_event)
		ni0O1li <= 1;
	always @(ni0O1ll_event)
		ni0O1ll <= 1;
	always @(ni0O1lO_event)
		ni0O1lO <= 1;
	always @(ni0O1Oi_event)
		ni0O1Oi <= 1;
	always @(ni0O1Ol_event)
		ni0O1Ol <= 1;
	always @(ni0O1OO_event)
		ni0O1OO <= 1;
	always @(ni0Oi0l_event)
		ni0Oi0l <= 1;
	always @(ni0Oi1i_event)
		ni0Oi1i <= 1;
	always @(ni0Oi1l_event)
		ni0Oi1l <= 1;
	always @(nii110i_event)
		nii110i <= 1;
	initial
	begin
		nii100i = 0;
		nii100l = 0;
		nii100O = 0;
		nii101i = 0;
		nii101l = 0;
		nii101O = 0;
		nii10ii = 0;
		nii10il = 0;
		nii10iO = 0;
		nii10li = 0;
		nii10ll = 0;
		nii10lO = 0;
		nii10Oi = 0;
		nii10Ol = 0;
		nii10OO = 0;
		nii11lO = 0;
		nii11Oi = 0;
		nii11Ol = 0;
		nii11OO = 0;
		nii1i0i = 0;
		nii1i0l = 0;
		nii1i1i = 0;
		nii1i1l = 0;
		nii1i1O = 0;
		nii1iii = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nii100i <= 0;
			nii100l <= 0;
			nii100O <= 0;
			nii101i <= 0;
			nii101l <= 0;
			nii101O <= 0;
			nii10ii <= 0;
			nii10il <= 0;
			nii10iO <= 0;
			nii10li <= 0;
			nii10ll <= 0;
			nii10lO <= 0;
			nii10Oi <= 0;
			nii10Ol <= 0;
			nii10OO <= 0;
			nii11lO <= 0;
			nii11Oi <= 0;
			nii11Ol <= 0;
			nii11OO <= 0;
			nii1i0i <= 0;
			nii1i0l <= 0;
			nii1i1i <= 0;
			nii1i1l <= 0;
			nii1i1O <= 0;
			nii1iii <= 0;
		end
		else if  (n0OOOOl == 1'b1) 
		begin
			nii100i <= ni0O1OO;
			nii100l <= ni0O01i;
			nii100O <= ni0O01l;
			nii101i <= ni0O1lO;
			nii101l <= ni0O1Oi;
			nii101O <= ni0O1Ol;
			nii10ii <= ni0O01O;
			nii10il <= ni0O00i;
			nii10iO <= ni0O00l;
			nii10li <= ni0O00O;
			nii10ll <= ni0O0ii;
			nii10lO <= ni0O0il;
			nii10Oi <= ni0O0iO;
			nii10Ol <= ni0O0li;
			nii10OO <= ni0O0ll;
			nii11lO <= nii110i;
			nii11Oi <= ni0O1iO;
			nii11Ol <= ni0O1li;
			nii11OO <= ni0O1ll;
			nii1i0i <= ni0O0OO;
			nii1i0l <= ni0Oi1i;
			nii1i1i <= ni0O0lO;
			nii1i1l <= ni0O0Oi;
			nii1i1O <= ni0O0Ol;
			nii1iii <= ni0Oi1l;
		end
	end
	event nii100i_event;
	event nii100l_event;
	event nii100O_event;
	event nii101i_event;
	event nii101l_event;
	event nii101O_event;
	event nii10ii_event;
	event nii10il_event;
	event nii10iO_event;
	event nii10li_event;
	event nii10ll_event;
	event nii10lO_event;
	event nii10Oi_event;
	event nii10Ol_event;
	event nii10OO_event;
	event nii11lO_event;
	event nii11Oi_event;
	event nii11Ol_event;
	event nii11OO_event;
	event nii1i0i_event;
	event nii1i0l_event;
	event nii1i1i_event;
	event nii1i1l_event;
	event nii1i1O_event;
	event nii1iii_event;
	initial
		#1 ->nii100i_event;
	initial
		#1 ->nii100l_event;
	initial
		#1 ->nii100O_event;
	initial
		#1 ->nii101i_event;
	initial
		#1 ->nii101l_event;
	initial
		#1 ->nii101O_event;
	initial
		#1 ->nii10ii_event;
	initial
		#1 ->nii10il_event;
	initial
		#1 ->nii10iO_event;
	initial
		#1 ->nii10li_event;
	initial
		#1 ->nii10ll_event;
	initial
		#1 ->nii10lO_event;
	initial
		#1 ->nii10Oi_event;
	initial
		#1 ->nii10Ol_event;
	initial
		#1 ->nii10OO_event;
	initial
		#1 ->nii11lO_event;
	initial
		#1 ->nii11Oi_event;
	initial
		#1 ->nii11Ol_event;
	initial
		#1 ->nii11OO_event;
	initial
		#1 ->nii1i0i_event;
	initial
		#1 ->nii1i0l_event;
	initial
		#1 ->nii1i1i_event;
	initial
		#1 ->nii1i1l_event;
	initial
		#1 ->nii1i1O_event;
	initial
		#1 ->nii1iii_event;
	always @(nii100i_event)
		nii100i <= 1;
	always @(nii100l_event)
		nii100l <= 1;
	always @(nii100O_event)
		nii100O <= 1;
	always @(nii101i_event)
		nii101i <= 1;
	always @(nii101l_event)
		nii101l <= 1;
	always @(nii101O_event)
		nii101O <= 1;
	always @(nii10ii_event)
		nii10ii <= 1;
	always @(nii10il_event)
		nii10il <= 1;
	always @(nii10iO_event)
		nii10iO <= 1;
	always @(nii10li_event)
		nii10li <= 1;
	always @(nii10ll_event)
		nii10ll <= 1;
	always @(nii10lO_event)
		nii10lO <= 1;
	always @(nii10Oi_event)
		nii10Oi <= 1;
	always @(nii10Ol_event)
		nii10Ol <= 1;
	always @(nii10OO_event)
		nii10OO <= 1;
	always @(nii11lO_event)
		nii11lO <= 1;
	always @(nii11Oi_event)
		nii11Oi <= 1;
	always @(nii11Ol_event)
		nii11Ol <= 1;
	always @(nii11OO_event)
		nii11OO <= 1;
	always @(nii1i0i_event)
		nii1i0i <= 1;
	always @(nii1i0l_event)
		nii1i0l <= 1;
	always @(nii1i1i_event)
		nii1i1i <= 1;
	always @(nii1i1l_event)
		nii1i1l <= 1;
	always @(nii1i1O_event)
		nii1i1O <= 1;
	always @(nii1iii_event)
		nii1iii <= 1;
	initial
	begin
		nii1iiO = 0;
		nii1ili = 0;
		nii1ill = 0;
		nii1ilO = 0;
		nii1iOi = 0;
		nii1iOl = 0;
		nii1iOO = 0;
		nii1l0i = 0;
		nii1l1i = 0;
		nii1l1l = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nii1iiO <= 0;
			nii1ili <= 0;
			nii1ill <= 0;
			nii1ilO <= 0;
			nii1iOi <= 0;
			nii1iOl <= 0;
			nii1iOO <= 0;
			nii1l0i <= 0;
			nii1l1i <= 0;
			nii1l1l <= 0;
		end
		else if  (n0OOOOO == 1'b1) 
		begin
			nii1iiO <= nl01i1i;
			nii1ili <= nl01i1l;
			nii1ill <= nl01i1O;
			nii1ilO <= nl01i0l;
			nii1iOi <= nl0101l;
			nii1iOl <= nl0101O;
			nii1iOO <= nl0100i;
			nii1l0i <= nl011ii;
			nii1l1i <= nl0100O;
			nii1l1l <= nl0110l;
		end
	end
	initial
	begin
		nii1lii = 0;
		nii1lil = 0;
		nii1liO = 0;
		nii1lli = 0;
		nii1lll = 0;
		nii1llO = 0;
		nii1lOi = 0;
		nii1lOO = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nii1lii <= 0;
			nii1lil <= 0;
			nii1liO <= 0;
			nii1lli <= 0;
			nii1lll <= 0;
			nii1llO <= 0;
			nii1lOi <= 0;
			nii1lOO <= 0;
		end
		else if  (ni1111i == 1'b1) 
		begin
			nii1lii <= nl01i1i;
			nii1lil <= nl01i1l;
			nii1liO <= nl01i1O;
			nii1lli <= nl01i0l;
			nii1lll <= nl0101l;
			nii1llO <= nl0101O;
			nii1lOi <= nl0100i;
			nii1lOO <= nl0100O;
		end
	end
	initial
	begin
		nii1O0i = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nii1O0i <= 0;
		end
		else if  (wire_nii1O1O_ENA == 1'b1) 
		begin
			nii1O0i <= nii1iii;
		end
	end
	assign
		wire_nii1O1O_ENA = (nlOOOl & (~ ni1iiii));
	initial
	begin
		nii1Oil = 0;
		nii1OiO = 0;
		nii1Oli = 0;
		nii1OlO = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nii1Oil <= 0;
			nii1OiO <= 0;
			nii1Oli <= 0;
			nii1OlO <= 0;
		end
		else if  (ni1111l == 1'b1) 
		begin
			nii1Oil <= wire_nii1OOl_dataout;
			nii1OiO <= wire_nii1OOO_dataout;
			nii1Oli <= wire_nii011i_dataout;
			nii1OlO <= wire_nii1OOi_dataout;
		end
	end
	initial
	begin
		nil10lO = 0;
		nil1i0i = 0;
		nil1i0l = 0;
		nil1i0O = 0;
		nil1i1O = 0;
		nil1iii = 0;
		nil1iil = 0;
		nil1iiO = 0;
		nil1ili = 0;
		nil1ill = 0;
		nil1ilO = 0;
		nil1iOi = 0;
		nil1iOl = 0;
		nil1iOO = 0;
		nil1l0i = 0;
		nil1l0l = 0;
		nil1l0O = 0;
		nil1l1i = 0;
		nil1l1l = 0;
		nil1l1O = 0;
		nil1lii = 0;
		nil1lil = 0;
		nil1liO = 0;
		nil1lli = 0;
		nil1llO = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nil10lO <= 0;
			nil1i0i <= 0;
			nil1i0l <= 0;
			nil1i0O <= 0;
			nil1i1O <= 0;
			nil1iii <= 0;
			nil1iil <= 0;
			nil1iiO <= 0;
			nil1ili <= 0;
			nil1ill <= 0;
			nil1ilO <= 0;
			nil1iOi <= 0;
			nil1iOl <= 0;
			nil1iOO <= 0;
			nil1l0i <= 0;
			nil1l0l <= 0;
			nil1l0O <= 0;
			nil1l1i <= 0;
			nil1l1l <= 0;
			nil1l1O <= 0;
			nil1lii <= 0;
			nil1lil <= 0;
			nil1liO <= 0;
			nil1lli <= 0;
			nil1llO <= 0;
		end
		else if  (ni110ii == 1'b1) 
		begin
			nil10lO <= wire_nilllii_dataout;
			nil1i0i <= wire_nill0Ol_dataout;
			nil1i0l <= wire_nill0OO_dataout;
			nil1i0O <= wire_nilli1i_dataout;
			nil1i1O <= wire_nill0Oi_dataout;
			nil1iii <= wire_nilli1l_dataout;
			nil1iil <= wire_nilli1O_dataout;
			nil1iiO <= wire_nilli0i_dataout;
			nil1ili <= wire_nilli0l_dataout;
			nil1ill <= wire_nilli0O_dataout;
			nil1ilO <= wire_nilliii_dataout;
			nil1iOi <= wire_nilliil_dataout;
			nil1iOl <= wire_nilliiO_dataout;
			nil1iOO <= wire_nillili_dataout;
			nil1l0i <= wire_nilliOl_dataout;
			nil1l0l <= wire_nilliOO_dataout;
			nil1l0O <= wire_nilll1i_dataout;
			nil1l1i <= wire_nillill_dataout;
			nil1l1l <= wire_nillilO_dataout;
			nil1l1O <= wire_nilliOi_dataout;
			nil1lii <= wire_nilll1l_dataout;
			nil1lil <= wire_nilll1O_dataout;
			nil1liO <= wire_nilll0i_dataout;
			nil1lli <= wire_nilll0l_dataout;
			nil1llO <= wire_nilll0O_dataout;
		end
	end
	event nil10lO_event;
	event nil1i0i_event;
	event nil1i0l_event;
	event nil1i0O_event;
	event nil1i1O_event;
	event nil1iii_event;
	event nil1iil_event;
	event nil1iiO_event;
	event nil1ili_event;
	event nil1ill_event;
	event nil1ilO_event;
	event nil1iOi_event;
	event nil1iOl_event;
	event nil1iOO_event;
	event nil1l0i_event;
	event nil1l0l_event;
	event nil1l0O_event;
	event nil1l1i_event;
	event nil1l1l_event;
	event nil1l1O_event;
	event nil1lii_event;
	event nil1lil_event;
	event nil1liO_event;
	event nil1lli_event;
	event nil1llO_event;
	initial
		#1 ->nil10lO_event;
	initial
		#1 ->nil1i0i_event;
	initial
		#1 ->nil1i0l_event;
	initial
		#1 ->nil1i0O_event;
	initial
		#1 ->nil1i1O_event;
	initial
		#1 ->nil1iii_event;
	initial
		#1 ->nil1iil_event;
	initial
		#1 ->nil1iiO_event;
	initial
		#1 ->nil1ili_event;
	initial
		#1 ->nil1ill_event;
	initial
		#1 ->nil1ilO_event;
	initial
		#1 ->nil1iOi_event;
	initial
		#1 ->nil1iOl_event;
	initial
		#1 ->nil1iOO_event;
	initial
		#1 ->nil1l0i_event;
	initial
		#1 ->nil1l0l_event;
	initial
		#1 ->nil1l0O_event;
	initial
		#1 ->nil1l1i_event;
	initial
		#1 ->nil1l1l_event;
	initial
		#1 ->nil1l1O_event;
	initial
		#1 ->nil1lii_event;
	initial
		#1 ->nil1lil_event;
	initial
		#1 ->nil1liO_event;
	initial
		#1 ->nil1lli_event;
	initial
		#1 ->nil1llO_event;
	always @(nil10lO_event)
		nil10lO <= 1;
	always @(nil1i0i_event)
		nil1i0i <= 1;
	always @(nil1i0l_event)
		nil1i0l <= 1;
	always @(nil1i0O_event)
		nil1i0O <= 1;
	always @(nil1i1O_event)
		nil1i1O <= 1;
	always @(nil1iii_event)
		nil1iii <= 1;
	always @(nil1iil_event)
		nil1iil <= 1;
	always @(nil1iiO_event)
		nil1iiO <= 1;
	always @(nil1ili_event)
		nil1ili <= 1;
	always @(nil1ill_event)
		nil1ill <= 1;
	always @(nil1ilO_event)
		nil1ilO <= 1;
	always @(nil1iOi_event)
		nil1iOi <= 1;
	always @(nil1iOl_event)
		nil1iOl <= 1;
	always @(nil1iOO_event)
		nil1iOO <= 1;
	always @(nil1l0i_event)
		nil1l0i <= 1;
	always @(nil1l0l_event)
		nil1l0l <= 1;
	always @(nil1l0O_event)
		nil1l0O <= 1;
	always @(nil1l1i_event)
		nil1l1i <= 1;
	always @(nil1l1l_event)
		nil1l1l <= 1;
	always @(nil1l1O_event)
		nil1l1O <= 1;
	always @(nil1lii_event)
		nil1lii <= 1;
	always @(nil1lil_event)
		nil1lil <= 1;
	always @(nil1liO_event)
		nil1liO <= 1;
	always @(nil1lli_event)
		nil1lli <= 1;
	always @(nil1llO_event)
		nil1llO <= 1;
	initial
	begin
		nilOiOl = 0;
		nilOl0l = 0;
		nilOl0O = 0;
		nilOlii = 0;
		nilOlil = 0;
		nilOliO = 0;
		nilOlli = 0;
		nilOlll = 0;
		nilOlOi = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nilOiOl <= 0;
			nilOl0l <= 0;
			nilOl0O <= 0;
			nilOlii <= 0;
			nilOlil <= 0;
			nilOliO <= 0;
			nilOlli <= 0;
			nilOlll <= 0;
			nilOlOi <= 0;
		end
		else if  (ni11iii == 1'b1) 
		begin
			nilOiOl <= wire_niO1OOO_dataout;
			nilOl0l <= wire_niO1Oii_dataout;
			nilOl0O <= wire_niO1Oil_dataout;
			nilOlii <= wire_niO1OiO_dataout;
			nilOlil <= wire_niO1Oli_dataout;
			nilOliO <= wire_niO1Oll_dataout;
			nilOlli <= wire_niO1OlO_dataout;
			nilOlll <= wire_niO1OOi_dataout;
			nilOlOi <= wire_niO1OOl_dataout;
		end
	end
	initial
	begin
		niOii1l = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			niOii1l <= 0;
		end
		else if  (wire_niOii1i_ENA == 1'b1) 
		begin
			niOii1l <= wire_niOi0Oi_o;
		end
	end
	assign
		wire_niOii1i_ENA = (wire_niOi00O_o & ni1iiiO);
	event niOii1l_event;
	initial
		#1 ->niOii1l_event;
	always @(niOii1l_event)
		niOii1l <= 1;
	initial
	begin
		niOii0i = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			niOii0i <= 1;
		end
		else if  (niOiOii == 1'b1) 
		begin
			niOii0i <= niOii1l;
		end
	end
	event niOii0i_event;
	initial
		#1 ->niOii0i_event;
	always @(niOii0i_event)
		niOii0i <= 1;
	initial
	begin
		niOiill = 0;
		niOiilO = 0;
		niOiiOi = 0;
		niOiiOl = 0;
		niOiiOO = 0;
		niOil0i = 0;
		niOil0l = 0;
		niOil0O = 0;
		niOil1i = 0;
		niOil1l = 0;
		niOil1O = 0;
		niOilii = 0;
		niOilil = 0;
		niOiliO = 0;
		niOilli = 0;
		niOilll = 0;
		niOillO = 0;
		niOilOi = 0;
		niOilOl = 0;
		niOilOO = 0;
		niOiO0l = 0;
		niOiO1i = 0;
		niOiO1l = 0;
		niOiO1O = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			niOiill <= 0;
			niOiilO <= 0;
			niOiiOi <= 0;
			niOiiOl <= 0;
			niOiiOO <= 0;
			niOil0i <= 0;
			niOil0l <= 0;
			niOil0O <= 0;
			niOil1i <= 0;
			niOil1l <= 0;
			niOil1O <= 0;
			niOilii <= 0;
			niOilil <= 0;
			niOiliO <= 0;
			niOilli <= 0;
			niOilll <= 0;
			niOillO <= 0;
			niOilOi <= 0;
			niOilOl <= 0;
			niOilOO <= 0;
			niOiO0l <= 0;
			niOiO1i <= 0;
			niOiO1l <= 0;
			niOiO1O <= 0;
		end
		else if  (ni11O0O == 1'b1) 
		begin
			niOiill <= wire_niO0O0O_o;
			niOiilO <= wire_niO0Oii_o;
			niOiiOi <= wire_niO0Oil_o;
			niOiiOl <= wire_niO0OiO_o;
			niOiiOO <= wire_niO0Oli_o;
			niOil0i <= wire_niO0OOl_o;
			niOil0l <= wire_niO0OOO_o;
			niOil0O <= wire_niOi11i_o;
			niOil1i <= wire_niO0Oll_o;
			niOil1l <= wire_niO0OlO_o;
			niOil1O <= wire_niO0OOi_o;
			niOilii <= wire_niOi11l_o;
			niOilil <= wire_niOi11O_o;
			niOiliO <= wire_niOi10i_o;
			niOilli <= wire_niOi10l_o;
			niOilll <= wire_niOi10O_o;
			niOillO <= wire_niOi1ii_o;
			niOilOi <= wire_niOi1il_o;
			niOilOl <= wire_niOi1iO_o;
			niOilOO <= wire_niOi1li_o;
			niOiO0l <= wire_niOi1Ol_o;
			niOiO1i <= wire_niOi1ll_o;
			niOiO1l <= wire_niOi1lO_o;
			niOiO1O <= wire_niOi1Oi_o;
		end
	end
	event niOiill_event;
	event niOiilO_event;
	event niOiiOi_event;
	event niOiiOl_event;
	event niOiiOO_event;
	event niOil0i_event;
	event niOil0l_event;
	event niOil0O_event;
	event niOil1i_event;
	event niOil1l_event;
	event niOil1O_event;
	event niOilii_event;
	event niOilil_event;
	event niOiliO_event;
	event niOilli_event;
	event niOilll_event;
	event niOillO_event;
	event niOilOi_event;
	event niOilOl_event;
	event niOilOO_event;
	event niOiO0l_event;
	event niOiO1i_event;
	event niOiO1l_event;
	event niOiO1O_event;
	initial
		#1 ->niOiill_event;
	initial
		#1 ->niOiilO_event;
	initial
		#1 ->niOiiOi_event;
	initial
		#1 ->niOiiOl_event;
	initial
		#1 ->niOiiOO_event;
	initial
		#1 ->niOil0i_event;
	initial
		#1 ->niOil0l_event;
	initial
		#1 ->niOil0O_event;
	initial
		#1 ->niOil1i_event;
	initial
		#1 ->niOil1l_event;
	initial
		#1 ->niOil1O_event;
	initial
		#1 ->niOilii_event;
	initial
		#1 ->niOilil_event;
	initial
		#1 ->niOiliO_event;
	initial
		#1 ->niOilli_event;
	initial
		#1 ->niOilll_event;
	initial
		#1 ->niOillO_event;
	initial
		#1 ->niOilOi_event;
	initial
		#1 ->niOilOl_event;
	initial
		#1 ->niOilOO_event;
	initial
		#1 ->niOiO0l_event;
	initial
		#1 ->niOiO1i_event;
	initial
		#1 ->niOiO1l_event;
	initial
		#1 ->niOiO1O_event;
	always @(niOiill_event)
		niOiill <= 1;
	always @(niOiilO_event)
		niOiilO <= 1;
	always @(niOiiOi_event)
		niOiiOi <= 1;
	always @(niOiiOl_event)
		niOiiOl <= 1;
	always @(niOiiOO_event)
		niOiiOO <= 1;
	always @(niOil0i_event)
		niOil0i <= 1;
	always @(niOil0l_event)
		niOil0l <= 1;
	always @(niOil0O_event)
		niOil0O <= 1;
	always @(niOil1i_event)
		niOil1i <= 1;
	always @(niOil1l_event)
		niOil1l <= 1;
	always @(niOil1O_event)
		niOil1O <= 1;
	always @(niOilii_event)
		niOilii <= 1;
	always @(niOilil_event)
		niOilil <= 1;
	always @(niOiliO_event)
		niOiliO <= 1;
	always @(niOilli_event)
		niOilli <= 1;
	always @(niOilll_event)
		niOilll <= 1;
	always @(niOillO_event)
		niOillO <= 1;
	always @(niOilOi_event)
		niOilOi <= 1;
	always @(niOilOl_event)
		niOilOl <= 1;
	always @(niOilOO_event)
		niOilOO <= 1;
	always @(niOiO0l_event)
		niOiO0l <= 1;
	always @(niOiO1i_event)
		niOiO1i <= 1;
	always @(niOiO1l_event)
		niOiO1l <= 1;
	always @(niOiO1O_event)
		niOiO1O <= 1;
	initial
	begin
		ni0000l = 0;
		ni0001i = 0;
		ni0001O = 0;
		ni000il = 0;
		ni000li = 0;
		ni000lO = 0;
		ni0011l = 0;
		ni001ii = 0;
		ni001ll = 0;
		ni001Ol = 0;
		ni00i0O = 0;
		ni00i1l = 0;
		ni00iiO = 0;
		ni00ill = 0;
		ni00iOi = 0;
		ni00iOO = 0;
		ni00l0l = 0;
		ni00l1O = 0;
		ni00lii = 0;
		ni00llO = 0;
		ni00O0i = 0;
		ni00O0O = 0;
		ni00O1i = 0;
		ni00Oil = 0;
		ni0100l = 0;
		ni010ii = 0;
		ni01i1O = 0;
		ni01iii = 0;
		ni01iil = 0;
		ni01liO = 0;
		ni01lli = 0;
		ni01Oli = 0;
		ni01OOi = 0;
		ni01OOO = 0;
		ni0Oi0i = 0;
		ni0Oi1O = 0;
		nii0lll = 0;
		nii0lOi = 0;
		nii0lOl = 0;
		nii0lOO = 0;
		nii0O0i = 0;
		nii0O0l = 0;
		nii0O0O = 0;
		nii0O1i = 0;
		nii0O1l = 0;
		nii0O1O = 0;
		nii0Oii = 0;
		nii0Oil = 0;
		nii0OiO = 0;
		nii0Oli = 0;
		nii0Oll = 0;
		nii0OlO = 0;
		nii0OOi = 0;
		nii0OOl = 0;
		nii0OOO = 0;
		niii00i = 0;
		niii00l = 0;
		niii00O = 0;
		niii01i = 0;
		niii01l = 0;
		niii01O = 0;
		niii0ii = 0;
		niii0il = 0;
		niii0iO = 0;
		niii0li = 0;
		niii0ll = 0;
		niii0lO = 0;
		niii0Oi = 0;
		niii0Ol = 0;
		niii0OO = 0;
		niii10i = 0;
		niii10l = 0;
		niii10O = 0;
		niii11i = 0;
		niii11l = 0;
		niii11O = 0;
		niii1ii = 0;
		niii1il = 0;
		niii1iO = 0;
		niii1li = 0;
		niii1ll = 0;
		niii1lO = 0;
		niii1Oi = 0;
		niii1Ol = 0;
		niii1OO = 0;
		niiii0i = 0;
		niiii0l = 0;
		niiii0O = 0;
		niiii1i = 0;
		niiii1l = 0;
		niiii1O = 0;
		niiiiii = 0;
		niiiiil = 0;
		niiiiiO = 0;
		niiiili = 0;
		niiiill = 0;
		niiiilO = 0;
		niiiiOi = 0;
		niiiiOl = 0;
		niiiiOO = 0;
		niiil0i = 0;
		niiil0l = 0;
		niiil0O = 0;
		niiil1i = 0;
		niiil1l = 0;
		niiil1O = 0;
		niiilii = 0;
		niiilil = 0;
		niiiliO = 0;
		niiilli = 0;
		niiilll = 0;
		niiillO = 0;
		niiilOi = 0;
		niiilOl = 0;
		nil000i = 0;
		nil000l = 0;
		nil000O = 0;
		nil001i = 0;
		nil001l = 0;
		nil001O = 0;
		nil00ii = 0;
		nil00il = 0;
		nil00iO = 0;
		nil00li = 0;
		nil00ll = 0;
		nil00lO = 0;
		nil00Oi = 0;
		nil00Ol = 0;
		nil00OO = 0;
		nil010i = 0;
		nil010l = 0;
		nil010O = 0;
		nil011i = 0;
		nil011l = 0;
		nil011O = 0;
		nil01ii = 0;
		nil01il = 0;
		nil01iO = 0;
		nil01li = 0;
		nil01ll = 0;
		nil01lO = 0;
		nil01Oi = 0;
		nil01Ol = 0;
		nil01OO = 0;
		nil0i0i = 0;
		nil0i0l = 0;
		nil0i0O = 0;
		nil0i1i = 0;
		nil0i1l = 0;
		nil0i1O = 0;
		nil0iii = 0;
		nil0iil = 0;
		nil0iiO = 0;
		nil0ili = 0;
		nil0ill = 0;
		nil0ilO = 0;
		nil0iOi = 0;
		nil0iOl = 0;
		nil0iOO = 0;
		nil0l0i = 0;
		nil0l0l = 0;
		nil0l0O = 0;
		nil0l1i = 0;
		nil0l1l = 0;
		nil0l1O = 0;
		nil0lii = 0;
		nil0lil = 0;
		nil0liO = 0;
		nil0lli = 0;
		nil0lll = 0;
		nil0llO = 0;
		nil0lOi = 0;
		nil0lOl = 0;
		nil0lOO = 0;
		nil0O1i = 0;
		nil101O = 0;
		nil11Ol = 0;
		nil11OO = 0;
		nil1lOi = 0;
		nil1lOO = 0;
		nil1O0i = 0;
		nil1O0l = 0;
		nil1O0O = 0;
		nil1O1i = 0;
		nil1O1l = 0;
		nil1O1O = 0;
		nil1Oii = 0;
		nil1Oil = 0;
		nil1OiO = 0;
		nil1Oli = 0;
		nil1Oll = 0;
		nil1OlO = 0;
		nil1OOi = 0;
		nil1OOl = 0;
		nil1OOO = 0;
		nilO00l = 0;
		nilO01i = 0;
		nilO01l = 0;
		nilO0iO = 0;
		nilO0li = 0;
		nilO0ll = 0;
		nilOi0l = 0;
		nilOlOl = 0;
		nilOO0i = 0;
		nilOO0l = 0;
		nilOO0O = 0;
		nilOO1i = 0;
		nilOO1l = 0;
		nilOO1O = 0;
		nilOOii = 0;
		nilOOil = 0;
		nilOOiO = 0;
		nilOOli = 0;
		nilOOll = 0;
		nilOOlO = 0;
		nilOOOi = 0;
		nilOOOl = 0;
		nilOOOO = 0;
		niO00il = 0;
		niO00iO = 0;
		niO00lO = 0;
		niO110i = 0;
		niO110l = 0;
		niO110O = 0;
		niO111i = 0;
		niO111l = 0;
		niO111O = 0;
		niO11ii = 0;
		niO11il = 0;
		niO11iO = 0;
		niO11li = 0;
		niO11ll = 0;
		niO11lO = 0;
		niO11Oi = 0;
		niO11Ol = 0;
		niOii0l = 0;
		niOiOii = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			ni0000l <= 0;
			ni0001i <= 0;
			ni0001O <= 0;
			ni000il <= 0;
			ni000li <= 0;
			ni000lO <= 0;
			ni0011l <= 0;
			ni001ii <= 0;
			ni001ll <= 0;
			ni001Ol <= 0;
			ni00i0O <= 0;
			ni00i1l <= 0;
			ni00iiO <= 0;
			ni00ill <= 0;
			ni00iOi <= 0;
			ni00iOO <= 0;
			ni00l0l <= 0;
			ni00l1O <= 0;
			ni00lii <= 0;
			ni00llO <= 0;
			ni00O0i <= 0;
			ni00O0O <= 0;
			ni00O1i <= 0;
			ni00Oil <= 0;
			ni0100l <= 0;
			ni010ii <= 0;
			ni01i1O <= 0;
			ni01iii <= 0;
			ni01iil <= 0;
			ni01liO <= 0;
			ni01lli <= 0;
			ni01Oli <= 0;
			ni01OOi <= 0;
			ni01OOO <= 0;
			ni0Oi0i <= 0;
			ni0Oi1O <= 0;
			nii0lll <= 0;
			nii0lOi <= 0;
			nii0lOl <= 0;
			nii0lOO <= 0;
			nii0O0i <= 0;
			nii0O0l <= 0;
			nii0O0O <= 0;
			nii0O1i <= 0;
			nii0O1l <= 0;
			nii0O1O <= 0;
			nii0Oii <= 0;
			nii0Oil <= 0;
			nii0OiO <= 0;
			nii0Oli <= 0;
			nii0Oll <= 0;
			nii0OlO <= 0;
			nii0OOi <= 0;
			nii0OOl <= 0;
			nii0OOO <= 0;
			niii00i <= 0;
			niii00l <= 0;
			niii00O <= 0;
			niii01i <= 0;
			niii01l <= 0;
			niii01O <= 0;
			niii0ii <= 0;
			niii0il <= 0;
			niii0iO <= 0;
			niii0li <= 0;
			niii0ll <= 0;
			niii0lO <= 0;
			niii0Oi <= 0;
			niii0Ol <= 0;
			niii0OO <= 0;
			niii10i <= 0;
			niii10l <= 0;
			niii10O <= 0;
			niii11i <= 0;
			niii11l <= 0;
			niii11O <= 0;
			niii1ii <= 0;
			niii1il <= 0;
			niii1iO <= 0;
			niii1li <= 0;
			niii1ll <= 0;
			niii1lO <= 0;
			niii1Oi <= 0;
			niii1Ol <= 0;
			niii1OO <= 0;
			niiii0i <= 0;
			niiii0l <= 0;
			niiii0O <= 0;
			niiii1i <= 0;
			niiii1l <= 0;
			niiii1O <= 0;
			niiiiii <= 0;
			niiiiil <= 0;
			niiiiiO <= 0;
			niiiili <= 0;
			niiiill <= 0;
			niiiilO <= 0;
			niiiiOi <= 0;
			niiiiOl <= 0;
			niiiiOO <= 0;
			niiil0i <= 0;
			niiil0l <= 0;
			niiil0O <= 0;
			niiil1i <= 0;
			niiil1l <= 0;
			niiil1O <= 0;
			niiilii <= 0;
			niiilil <= 0;
			niiiliO <= 0;
			niiilli <= 0;
			niiilll <= 0;
			niiillO <= 0;
			niiilOi <= 0;
			niiilOl <= 0;
			nil000i <= 0;
			nil000l <= 0;
			nil000O <= 0;
			nil001i <= 0;
			nil001l <= 0;
			nil001O <= 0;
			nil00ii <= 0;
			nil00il <= 0;
			nil00iO <= 0;
			nil00li <= 0;
			nil00ll <= 0;
			nil00lO <= 0;
			nil00Oi <= 0;
			nil00Ol <= 0;
			nil00OO <= 0;
			nil010i <= 0;
			nil010l <= 0;
			nil010O <= 0;
			nil011i <= 0;
			nil011l <= 0;
			nil011O <= 0;
			nil01ii <= 0;
			nil01il <= 0;
			nil01iO <= 0;
			nil01li <= 0;
			nil01ll <= 0;
			nil01lO <= 0;
			nil01Oi <= 0;
			nil01Ol <= 0;
			nil01OO <= 0;
			nil0i0i <= 0;
			nil0i0l <= 0;
			nil0i0O <= 0;
			nil0i1i <= 0;
			nil0i1l <= 0;
			nil0i1O <= 0;
			nil0iii <= 0;
			nil0iil <= 0;
			nil0iiO <= 0;
			nil0ili <= 0;
			nil0ill <= 0;
			nil0ilO <= 0;
			nil0iOi <= 0;
			nil0iOl <= 0;
			nil0iOO <= 0;
			nil0l0i <= 0;
			nil0l0l <= 0;
			nil0l0O <= 0;
			nil0l1i <= 0;
			nil0l1l <= 0;
			nil0l1O <= 0;
			nil0lii <= 0;
			nil0lil <= 0;
			nil0liO <= 0;
			nil0lli <= 0;
			nil0lll <= 0;
			nil0llO <= 0;
			nil0lOi <= 0;
			nil0lOl <= 0;
			nil0lOO <= 0;
			nil0O1i <= 0;
			nil101O <= 0;
			nil11Ol <= 0;
			nil11OO <= 0;
			nil1lOi <= 0;
			nil1lOO <= 0;
			nil1O0i <= 0;
			nil1O0l <= 0;
			nil1O0O <= 0;
			nil1O1i <= 0;
			nil1O1l <= 0;
			nil1O1O <= 0;
			nil1Oii <= 0;
			nil1Oil <= 0;
			nil1OiO <= 0;
			nil1Oli <= 0;
			nil1Oll <= 0;
			nil1OlO <= 0;
			nil1OOi <= 0;
			nil1OOl <= 0;
			nil1OOO <= 0;
			nilO00l <= 0;
			nilO01i <= 0;
			nilO01l <= 0;
			nilO0iO <= 0;
			nilO0li <= 0;
			nilO0ll <= 0;
			nilOi0l <= 0;
			nilOlOl <= 0;
			nilOO0i <= 0;
			nilOO0l <= 0;
			nilOO0O <= 0;
			nilOO1i <= 0;
			nilOO1l <= 0;
			nilOO1O <= 0;
			nilOOii <= 0;
			nilOOil <= 0;
			nilOOiO <= 0;
			nilOOli <= 0;
			nilOOll <= 0;
			nilOOlO <= 0;
			nilOOOi <= 0;
			nilOOOl <= 0;
			nilOOOO <= 0;
			niO00il <= 0;
			niO00iO <= 0;
			niO00lO <= 0;
			niO110i <= 0;
			niO110l <= 0;
			niO110O <= 0;
			niO111i <= 0;
			niO111l <= 0;
			niO111O <= 0;
			niO11ii <= 0;
			niO11il <= 0;
			niO11iO <= 0;
			niO11li <= 0;
			niO11ll <= 0;
			niO11lO <= 0;
			niO11Oi <= 0;
			niO11Ol <= 0;
			niOii0l <= 0;
			niOiOii <= 0;
		end
		else 
		begin
			ni0000l <= wire_ni0il0l_dataout;
			ni0001i <= wire_ni0ll0l_dataout;
			ni0001O <= wire_ni0llii_dataout;
			ni000il <= wire_ni0ilil_dataout;
			ni000li <= wire_ni0illi_dataout;
			ni000lO <= wire_ni0illO_dataout;
			ni0011l <= wire_ni0li0O_dataout;
			ni001ii <= wire_ni0lill_dataout;
			ni001ll <= wire_ni0liOO_dataout;
			ni001Ol <= wire_ni0ll1O_dataout;
			ni00i0O <= wire_ni0iO0O_dataout;
			ni00i1l <= wire_ni0iO1l_dataout;
			ni00iiO <= wire_ni0iOiO_dataout;
			ni00ill <= wire_ni0iOll_dataout;
			ni00iOi <= wire_ni0iOOi_dataout;
			ni00iOO <= wire_ni00Oli_dataout;
			ni00l0l <= wire_ni00OOO_dataout;
			ni00l1O <= wire_ni00OOi_dataout;
			ni00lii <= wire_ni0i11l_dataout;
			ni00llO <= wire_ni0i1ii_dataout;
			ni00O0i <= wire_ni0i1Ol_dataout;
			ni00O0O <= wire_ni0i01i_dataout;
			ni00O1i <= wire_ni0i1ll_dataout;
			ni00Oil <= wire_ni0i01O_dataout;
			ni0100l <= wire_ni010iO_dataout;
			ni010ii <= wire_ni01iiO_dataout;
			ni01i1O <= wire_ni010il_dataout;
			ni01iii <= wire_ni01ili_dataout;
			ni01iil <= wire_ni01iOi_dataout;
			ni01liO <= wire_ni01lll_dataout;
			ni01lli <= wire_ni01llO_dataout;
			ni01Oli <= wire_ni0l0Ol_dataout;
			ni01OOi <= wire_ni0li1l_dataout;
			ni01OOO <= wire_ni0li0i_dataout;
			ni0Oi0i <= wire_ni0O1il_dataout;
			ni0Oi1O <= wire_ni0Oi0O_dataout;
			nii0lll <= wire_niiO0iO_dataout;
			nii0lOi <= wire_niiliOi_dataout;
			nii0lOl <= wire_niiiO1i_dataout;
			nii0lOO <= wire_niiO0ll_dataout;
			nii0O0i <= wire_niiO0OO_dataout;
			nii0O0l <= wire_niiOi1i_dataout;
			nii0O0O <= wire_niiOi1l_dataout;
			nii0O1i <= wire_niiO0lO_dataout;
			nii0O1l <= wire_niiO0Oi_dataout;
			nii0O1O <= wire_niiO0Ol_dataout;
			nii0Oii <= wire_niiOi1O_dataout;
			nii0Oil <= wire_niiOi0i_dataout;
			nii0OiO <= wire_niiOi0l_dataout;
			nii0Oli <= wire_niiOi0O_dataout;
			nii0Oll <= wire_niiOiii_dataout;
			nii0OlO <= wire_niiOiil_dataout;
			nii0OOi <= wire_niiOiiO_dataout;
			nii0OOl <= wire_niiOili_dataout;
			nii0OOO <= wire_niiOill_dataout;
			niii00i <= wire_niilliO_dataout;
			niii00l <= wire_niillli_dataout;
			niii00O <= wire_niillll_dataout;
			niii01i <= wire_niill0O_dataout;
			niii01l <= wire_niillii_dataout;
			niii01O <= wire_niillil_dataout;
			niii0ii <= wire_niilllO_dataout;
			niii0il <= wire_niillOi_dataout;
			niii0iO <= wire_niillOl_dataout;
			niii0li <= wire_niillOO_dataout;
			niii0ll <= wire_niilO1i_dataout;
			niii0lO <= wire_niilO1l_dataout;
			niii0Oi <= wire_niilO1O_dataout;
			niii0Ol <= wire_niilO0i_dataout;
			niii0OO <= wire_niilO0l_dataout;
			niii10i <= wire_niiOiOO_dataout;
			niii10l <= wire_niiOl1i_dataout;
			niii10O <= wire_niiOl1l_dataout;
			niii11i <= wire_niiOilO_dataout;
			niii11l <= wire_niiOiOi_dataout;
			niii11O <= wire_niiOiOl_dataout;
			niii1ii <= wire_niiOl1O_dataout;
			niii1il <= wire_niiOl0i_dataout;
			niii1iO <= wire_niiOl0l_dataout;
			niii1li <= wire_niiliOO_dataout;
			niii1ll <= wire_niill1i_dataout;
			niii1lO <= wire_niill1l_dataout;
			niii1Oi <= wire_niill1O_dataout;
			niii1Ol <= wire_niill0i_dataout;
			niii1OO <= wire_niill0l_dataout;
			niiii0i <= wire_niilOiO_dataout;
			niiii0l <= wire_niiiO1O_dataout;
			niiii0O <= wire_niiiO0i_dataout;
			niiii1i <= wire_niilO0O_dataout;
			niiii1l <= wire_niilOii_dataout;
			niiii1O <= wire_niilOil_dataout;
			niiiiii <= wire_niiiO0l_dataout;
			niiiiil <= wire_niiiO0O_dataout;
			niiiiiO <= wire_niiiOii_dataout;
			niiiili <= wire_niiiOil_dataout;
			niiiill <= wire_niiiOiO_dataout;
			niiiilO <= wire_niiiOli_dataout;
			niiiiOi <= wire_niiiOll_dataout;
			niiiiOl <= wire_niiiOlO_dataout;
			niiiiOO <= wire_niiiOOi_dataout;
			niiil0i <= wire_niil11l_dataout;
			niiil0l <= wire_niil11O_dataout;
			niiil0O <= wire_niil10i_dataout;
			niiil1i <= wire_niiiOOl_dataout;
			niiil1l <= wire_niiiOOO_dataout;
			niiil1O <= wire_niil11i_dataout;
			niiilii <= wire_niil10l_dataout;
			niiilil <= wire_niil10O_dataout;
			niiiliO <= wire_niil1ii_dataout;
			niiilli <= wire_niil1il_dataout;
			niiilll <= wire_niil1iO_dataout;
			niiillO <= wire_niil1li_dataout;
			niiilOi <= wire_niil1ll_dataout;
			niiilOl <= wire_niil1lO_dataout;
			nil000i <= wire_nililiO_dataout;
			nil000l <= wire_nililli_dataout;
			nil000O <= wire_nililll_dataout;
			nil001i <= wire_nilil0O_dataout;
			nil001l <= wire_nililii_dataout;
			nil001O <= wire_nililil_dataout;
			nil00ii <= wire_nilillO_dataout;
			nil00il <= wire_nililOi_dataout;
			nil00iO <= wire_nililOl_dataout;
			nil00li <= wire_nililOO_dataout;
			nil00ll <= wire_niliO1i_dataout;
			nil00lO <= wire_niliO1l_dataout;
			nil00Oi <= wire_niliO1O_dataout;
			nil00Ol <= wire_niliO0i_dataout;
			nil00OO <= wire_niliO0l_dataout;
			nil010i <= wire_nilliOO_dataout;
			nil010l <= wire_nilll1i_dataout;
			nil010O <= wire_nilll1l_dataout;
			nil011i <= wire_nillilO_dataout;
			nil011l <= wire_nilliOi_dataout;
			nil011O <= wire_nilliOl_dataout;
			nil01ii <= wire_nilll1O_dataout;
			nil01il <= wire_nilll0i_dataout;
			nil01iO <= wire_nilll0l_dataout;
			nil01li <= wire_nilll0O_dataout;
			nil01ll <= wire_nilllii_dataout;
			nil01lO <= wire_nilil1l_dataout;
			nil01Oi <= wire_nilil1O_dataout;
			nil01Ol <= wire_nilil0i_dataout;
			nil01OO <= wire_nilil0l_dataout;
			nil0i0i <= wire_niliOiO_dataout;
			nil0i0l <= wire_niliOli_dataout;
			nil0i0O <= wire_niliOll_dataout;
			nil0i1i <= wire_niliO0O_dataout;
			nil0i1l <= wire_niliOii_dataout;
			nil0i1O <= wire_niliOil_dataout;
			nil0iii <= wire_nil0O0l_dataout;
			nil0iil <= wire_nil0O0O_dataout;
			nil0iiO <= wire_nil0Oii_dataout;
			nil0ili <= wire_nil0Oil_dataout;
			nil0ill <= wire_nil0OiO_dataout;
			nil0ilO <= wire_nil0Oli_dataout;
			nil0iOi <= wire_nil0Oll_dataout;
			nil0iOl <= wire_nil0OlO_dataout;
			nil0iOO <= wire_nil0OOi_dataout;
			nil0l0i <= wire_nili11l_dataout;
			nil0l0l <= wire_nili11O_dataout;
			nil0l0O <= wire_nili10i_dataout;
			nil0l1i <= wire_nil0OOl_dataout;
			nil0l1l <= wire_nil0OOO_dataout;
			nil0l1O <= wire_nili11i_dataout;
			nil0lii <= wire_nili10l_dataout;
			nil0lil <= wire_nili10O_dataout;
			nil0liO <= wire_nili1ii_dataout;
			nil0lli <= wire_nili1il_dataout;
			nil0lll <= wire_nili1iO_dataout;
			nil0llO <= wire_nili1li_dataout;
			nil0lOi <= wire_nili1ll_dataout;
			nil0lOl <= wire_nili1lO_dataout;
			nil0lOO <= wire_nili1Oi_dataout;
			nil0O1i <= wire_nili1Ol_dataout;
			nil101O <= wire_nii00ll_dataout;
			nil11Ol <= wire_nil101i_dataout;
			nil11OO <= wire_nil101l_dataout;
			nil1lOi <= wire_nill0ll_dataout;
			nil1lOO <= wire_niliiOO_dataout;
			nil1O0i <= wire_nill0OO_dataout;
			nil1O0l <= wire_nilli1i_dataout;
			nil1O0O <= wire_nilli1l_dataout;
			nil1O1i <= wire_nil0O1O_dataout;
			nil1O1l <= wire_nill0Oi_dataout;
			nil1O1O <= wire_nill0Ol_dataout;
			nil1Oii <= wire_nilli1O_dataout;
			nil1Oil <= wire_nilli0i_dataout;
			nil1OiO <= wire_nilli0l_dataout;
			nil1Oli <= wire_nilli0O_dataout;
			nil1Oll <= wire_nilliii_dataout;
			nil1OlO <= wire_nilliil_dataout;
			nil1OOi <= wire_nilliiO_dataout;
			nil1OOl <= wire_nillili_dataout;
			nil1OOO <= wire_nillill_dataout;
			nilO00l <= wire_nil10Oi_dataout;
			nilO01i <= wire_nilO01O_dataout;
			nilO01l <= wire_nilO00i_dataout;
			nilO0iO <= wire_nilOi1l_dataout;
			nilO0li <= wire_nilO0OO_dataout;
			nilO0ll <= wire_nilO0lO_dataout;
			nilOi0l <= wire_nilO00O_dataout;
			nilOlOl <= wire_niO1O0l_dataout;
			nilOO0i <= wire_niO1Oil_dataout;
			nilOO0l <= wire_niO1OiO_dataout;
			nilOO0O <= wire_niO1Oli_dataout;
			nilOO1i <= wire_niO1ill_dataout;
			nilOO1l <= wire_niO101i_dataout;
			nilOO1O <= wire_niO1Oii_dataout;
			nilOOii <= wire_niO1Oll_dataout;
			nilOOil <= wire_niO1OlO_dataout;
			nilOOiO <= wire_niO1OOi_dataout;
			nilOOli <= wire_niO1OOl_dataout;
			nilOOll <= wire_niO1OOO_dataout;
			nilOOlO <= wire_niO1iOi_dataout;
			nilOOOi <= wire_niO1iOl_dataout;
			nilOOOl <= wire_niO1iOO_dataout;
			nilOOOO <= wire_niO1l1i_dataout;
			niO00il <= wire_niO00li_dataout;
			niO00iO <= wire_niO00ll_dataout;
			niO00lO <= wire_nilOiOO_dataout;
			niO110i <= wire_niO1l0l_dataout;
			niO110l <= wire_niO1l0O_dataout;
			niO110O <= wire_niO101O_dataout;
			niO111i <= wire_niO1l1l_dataout;
			niO111l <= wire_niO1l1O_dataout;
			niO111O <= wire_niO1l0i_dataout;
			niO11ii <= wire_niO100i_dataout;
			niO11il <= wire_niO100l_dataout;
			niO11iO <= wire_niO100O_dataout;
			niO11li <= wire_niO10ii_dataout;
			niO11ll <= wire_niO10il_dataout;
			niO11lO <= wire_niO10iO_dataout;
			niO11Oi <= wire_niO10li_dataout;
			niO11Ol <= wire_niO10ll_dataout;
			niOii0l <= wire_niOiOil_dataout;
			niOiOii <= (dout_ready & (ni11Oii | niOii0l));
		end
	end
	initial
	begin
		niOl0Ol = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			niOl0Ol <= 0;
		end
		else if  (ni11Oll == 1'b1) 
		begin
			niOl0Ol <= n0Oii;
		end
	end
	initial
	begin
		niOl0OO = 0;
		niOli0i = 0;
		niOli0l = 0;
		niOli0O = 0;
		niOli1i = 0;
		niOli1l = 0;
		niOli1O = 0;
		niOliii = 0;
		niOliil = 0;
		niOlili = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			niOl0OO <= 0;
			niOli0i <= 0;
			niOli0l <= 0;
			niOli0O <= 0;
			niOli1i <= 0;
			niOli1l <= 0;
			niOli1O <= 0;
			niOliii <= 0;
			niOliil <= 0;
			niOlili <= 0;
		end
		else if  (ni11OlO == 1'b1) 
		begin
			niOl0OO <= wire_niOl0il_q_a[1];
			niOli0i <= wire_niOl0il_q_a[5];
			niOli0l <= wire_niOl0il_q_a[6];
			niOli0O <= wire_niOl0il_q_a[7];
			niOli1i <= wire_niOl0il_q_a[2];
			niOli1l <= wire_niOl0il_q_a[3];
			niOli1O <= wire_niOl0il_q_a[4];
			niOliii <= wire_niOl0il_q_a[8];
			niOliil <= wire_niOl0il_q_a[9];
			niOlili <= wire_niOl0il_q_a[0];
		end
	end
	initial
	begin
		niOlO0i = 0;
		niOlO0l = 0;
		niOlO0O = 0;
		niOlO1l = 0;
		niOlO1O = 0;
		niOlOii = 0;
		niOlOil = 0;
		niOlOiO = 0;
		niOlOli = 0;
		niOlOlO = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			niOlO0i <= 0;
			niOlO0l <= 0;
			niOlO0O <= 0;
			niOlO1l <= 0;
			niOlO1O <= 0;
			niOlOii <= 0;
			niOlOil <= 0;
			niOlOiO <= 0;
			niOlOli <= 0;
			niOlOlO <= 0;
		end
		else if  (ni11OOi == 1'b1) 
		begin
			niOlO0i <= wire_niOlliO_o;
			niOlO0l <= wire_niOllli_o;
			niOlO0O <= wire_niOllll_o;
			niOlO1l <= wire_niOllii_o;
			niOlO1O <= wire_niOllil_o;
			niOlOii <= wire_niOlllO_o;
			niOlOil <= wire_niOllOi_o;
			niOlOiO <= wire_niOllOl_o;
			niOlOli <= wire_niOllOO_o;
			niOlOlO <= wire_niOll0O_o;
		end
	end
	initial
	begin
		niOO00i = 0;
		niOO00l = 0;
		niOO01i = 0;
		niOO01l = 0;
		niOO01O = 0;
		niOO0ii = 0;
		niOO1Ol = 0;
		niOO1OO = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			niOO00i <= 0;
			niOO00l <= 0;
			niOO01i <= 0;
			niOO01l <= 0;
			niOO01O <= 0;
			niOO0ii <= 0;
			niOO1Ol <= 0;
			niOO1OO <= 0;
		end
		else if  (ni11OOO == 1'b1) 
		begin
			niOO00i <= wire_niOl0il_q_a[5];
			niOO00l <= wire_niOl0il_q_a[6];
			niOO01i <= wire_niOl0il_q_a[2];
			niOO01l <= wire_niOl0il_q_a[3];
			niOO01O <= wire_niOl0il_q_a[4];
			niOO0ii <= wire_niOl0il_q_a[7];
			niOO1Ol <= wire_niOl0il_q_a[0];
			niOO1OO <= wire_niOl0il_q_a[1];
		end
	end
	event niOO00i_event;
	event niOO00l_event;
	event niOO01i_event;
	event niOO01l_event;
	event niOO01O_event;
	event niOO0ii_event;
	event niOO1Ol_event;
	event niOO1OO_event;
	initial
		#1 ->niOO00i_event;
	initial
		#1 ->niOO00l_event;
	initial
		#1 ->niOO01i_event;
	initial
		#1 ->niOO01l_event;
	initial
		#1 ->niOO01O_event;
	initial
		#1 ->niOO0ii_event;
	initial
		#1 ->niOO1Ol_event;
	initial
		#1 ->niOO1OO_event;
	always @(niOO00i_event)
		niOO00i <= 1;
	always @(niOO00l_event)
		niOO00l <= 1;
	always @(niOO01i_event)
		niOO01i <= 1;
	always @(niOO01l_event)
		niOO01l <= 1;
	always @(niOO01O_event)
		niOO01O <= 1;
	always @(niOO0ii_event)
		niOO0ii <= 1;
	always @(niOO1Ol_event)
		niOO1Ol <= 1;
	always @(niOO1OO_event)
		niOO1OO <= 1;
	initial
	begin
		niOO10i = 0;
		niOO10l = 0;
		niOO10O = 0;
		niOO11i = 0;
		niOO11l = 0;
		niOO11O = 0;
		niOO1ii = 0;
		niOO1il = 0;
		niOO1iO = 0;
		niOO1ll = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			niOO10i <= 0;
			niOO10l <= 0;
			niOO10O <= 0;
			niOO11i <= 0;
			niOO11l <= 0;
			niOO11O <= 0;
			niOO1ii <= 0;
			niOO1il <= 0;
			niOO1iO <= 0;
			niOO1ll <= 0;
		end
		else if  (ni11OOl == 1'b1) 
		begin
			niOO10i <= wire_niOO1lO_o[5];
			niOO10l <= wire_niOO1lO_o[6];
			niOO10O <= wire_niOO1lO_o[7];
			niOO11i <= wire_niOO1lO_o[2];
			niOO11l <= wire_niOO1lO_o[3];
			niOO11O <= wire_niOO1lO_o[4];
			niOO1ii <= wire_niOO1lO_o[8];
			niOO1il <= wire_niOO1lO_o[9];
			niOO1iO <= wire_niOO1lO_o[10];
			niOO1ll <= wire_niOO1lO_o[1];
		end
	end
	initial
	begin
		niOO0ll = 0;
		niOO0lO = 0;
		niOO0Oi = 0;
		niOO0Ol = 0;
		niOO0OO = 0;
		niOOi0i = 0;
		niOOi1i = 0;
		niOOi1l = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			niOO0ll <= 0;
			niOO0lO <= 0;
			niOO0Oi <= 0;
			niOO0Ol <= 0;
			niOO0OO <= 0;
			niOOi0i <= 0;
			niOOi1i <= 0;
			niOOi1l <= 0;
		end
		else if  (ni1011i == 1'b1) 
		begin
			niOO0ll <= wire_niOOi0l_o[2];
			niOO0lO <= wire_niOOi0l_o[3];
			niOO0Oi <= wire_niOOi0l_o[4];
			niOO0Ol <= wire_niOOi0l_o[5];
			niOO0OO <= wire_niOOi0l_o[6];
			niOOi0i <= wire_niOOi0l_o[1];
			niOOi1i <= wire_niOOi0l_o[7];
			niOOi1l <= wire_niOOi0l_o[8];
		end
	end
	event niOO0ll_event;
	event niOO0lO_event;
	event niOO0Oi_event;
	event niOO0Ol_event;
	event niOO0OO_event;
	event niOOi0i_event;
	event niOOi1i_event;
	event niOOi1l_event;
	initial
		#1 ->niOO0ll_event;
	initial
		#1 ->niOO0lO_event;
	initial
		#1 ->niOO0Oi_event;
	initial
		#1 ->niOO0Ol_event;
	initial
		#1 ->niOO0OO_event;
	initial
		#1 ->niOOi0i_event;
	initial
		#1 ->niOOi1i_event;
	initial
		#1 ->niOOi1l_event;
	always @(niOO0ll_event)
		niOO0ll <= 1;
	always @(niOO0lO_event)
		niOO0lO <= 1;
	always @(niOO0Oi_event)
		niOO0Oi <= 1;
	always @(niOO0Ol_event)
		niOO0Ol <= 1;
	always @(niOO0OO_event)
		niOO0OO <= 1;
	always @(niOOi0i_event)
		niOOi0i <= 1;
	always @(niOOi1i_event)
		niOOi1i <= 1;
	always @(niOOi1l_event)
		niOOi1l <= 1;
	initial
	begin
		nl00i0l = 0;
		nl00i0O = 0;
		nl00iii = 0;
		nl00iil = 0;
		nl00iiO = 0;
		nl00ili = 0;
		nl00ill = 0;
		nl00ilO = 0;
		nl00iOi = 0;
		nl00iOO = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nl00i0l <= 0;
			nl00i0O <= 0;
			nl00iii <= 0;
			nl00iil <= 0;
			nl00iiO <= 0;
			nl00ili <= 0;
			nl00ill <= 0;
			nl00ilO <= 0;
			nl00iOi <= 0;
			nl00iOO <= 0;
		end
		else if  (ni10O1O == 1'b1) 
		begin
			nl00i0l <= wire_nl000iO_o;
			nl00i0O <= wire_nl000li_o;
			nl00iii <= wire_nl000ll_o;
			nl00iil <= wire_nl000lO_o;
			nl00iiO <= wire_nl000Oi_o;
			nl00ili <= wire_nl000Ol_o;
			nl00ill <= wire_nl000OO_o;
			nl00ilO <= wire_nl00i1i_o;
			nl00iOi <= wire_nl00i1l_o;
			nl00iOO <= wire_nl00i1O_o;
		end
	end
	initial
	begin
		nl00l0i = 0;
		nl00l0l = 0;
		nl00l0O = 0;
		nl00l1l = 0;
		nl00l1O = 0;
		nl00lil = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nl00l0i <= 0;
			nl00l0l <= 0;
			nl00l0O <= 0;
			nl00l1l <= 0;
			nl00l1O <= 0;
			nl00lil <= 0;
		end
		else if  (n0OiO == 1'b1) 
		begin
			nl00l0i <= nii010l;
			nl00l0l <= nii010O;
			nl00l0O <= nii01ii;
			nl00l1l <= nii01li;
			nl00l1O <= nii010i;
			nl00lil <= nii01il;
		end
	end
	event nl00l0i_event;
	event nl00l0l_event;
	event nl00l0O_event;
	event nl00l1l_event;
	event nl00l1O_event;
	event nl00lil_event;
	initial
		#1 ->nl00l0i_event;
	initial
		#1 ->nl00l0l_event;
	initial
		#1 ->nl00l0O_event;
	initial
		#1 ->nl00l1l_event;
	initial
		#1 ->nl00l1O_event;
	initial
		#1 ->nl00lil_event;
	always @(nl00l0i_event)
		nl00l0i <= 1;
	always @(nl00l0l_event)
		nl00l0l <= 1;
	always @(nl00l0O_event)
		nl00l0O <= 1;
	always @(nl00l1l_event)
		nl00l1l <= 1;
	always @(nl00l1O_event)
		nl00l1O <= 1;
	always @(nl00lil_event)
		nl00lil <= 1;
	initial
	begin
		nl00lli = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nl00lli <= 0;
		end
		else if  (wire_nl00liO_ENA == 1'b1) 
		begin
			nl00lli <= ni1il1i;
		end
	end
	assign
		wire_nl00liO_ENA = (n0Oll & (~ ni1iili));
	event nl00lli_event;
	initial
		#1 ->nl00lli_event;
	always @(nl00lli_event)
		nl00lli <= 1;
	initial
	begin
		nl00llO = 0;
		nl00lOi = 0;
		nl00lOl = 0;
		nl00O1i = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nl00llO <= 0;
			nl00lOi <= 0;
			nl00lOl <= 0;
			nl00O1i <= 0;
		end
		else if  (ni10O0i == 1'b1) 
		begin
			nl00llO <= nl1101l;
			nl00lOi <= nl1101O;
			nl00lOl <= nl1100i;
			nl00O1i <= nl1100l;
		end
	end
	initial
	begin
		nl00O0i = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nl00O0i <= 0;
		end
		else if  (wire_nl00O1O_ENA == 1'b1) 
		begin
			nl00O0i <= (nl1i0OO | nl1i0Oi);
		end
	end
	assign
		wire_nl00O1O_ENA = (n0Oll & (~ ni1iili));
	event nl00O0i_event;
	initial
		#1 ->nl00O0i_event;
	always @(nl00O0i_event)
		nl00O0i <= 1;
	initial
	begin
		nl00O0O = 0;
		nl00Oii = 0;
		nl00Oil = 0;
		nl00Oli = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nl00O0O <= 0;
			nl00Oii <= 0;
			nl00Oil <= 0;
			nl00Oli <= 0;
		end
		else if  (ni10O0l == 1'b1) 
		begin
			nl00O0O <= nl100iO;
			nl00Oii <= nl100li;
			nl00Oil <= nl100ll;
			nl00Oli <= nl100lO;
		end
	end
	initial
	begin
		nl0100i = 0;
		nl0100O = 0;
		nl0101l = 0;
		nl0101O = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nl0100i <= 0;
			nl0100O <= 0;
			nl0101l <= 0;
			nl0101O <= 0;
		end
		else if  (ni100lO == 1'b1) 
		begin
			nl0100i <= wire_nl011Ol_o;
			nl0100O <= wire_nl011OO_o;
			nl0101l <= wire_nl011lO_o;
			nl0101O <= wire_nl011Oi_o;
		end
	end
	event nl0100i_event;
	event nl0100O_event;
	event nl0101l_event;
	event nl0101O_event;
	initial
		#1 ->nl0100i_event;
	initial
		#1 ->nl0100O_event;
	initial
		#1 ->nl0101l_event;
	initial
		#1 ->nl0101O_event;
	always @(nl0100i_event)
		nl0100i <= 1;
	always @(nl0100O_event)
		nl0100O <= 1;
	always @(nl0101l_event)
		nl0101l <= 1;
	always @(nl0101O_event)
		nl0101O <= 1;
	initial
	begin
		nl0110l = 0;
		nl011ii = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nl0110l <= 0;
			nl011ii <= 0;
		end
		else if  (ni100ll == 1'b1) 
		begin
			nl0110l <= wire_nl0111l_o;
			nl011ii <= wire_nl0111O_o;
		end
	end
	event nl0110l_event;
	event nl011ii_event;
	initial
		#1 ->nl0110l_event;
	initial
		#1 ->nl011ii_event;
	always @(nl0110l_event)
		nl0110l <= 1;
	always @(nl011ii_event)
		nl011ii <= 1;
	initial
	begin
		nl01i0l = 0;
		nl01i1i = 0;
		nl01i1l = 0;
		nl01i1O = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nl01i0l <= 0;
			nl01i1i <= 0;
			nl01i1l <= 0;
			nl01i1O <= 0;
		end
		else if  (ni100Oi == 1'b1) 
		begin
			nl01i0l <= wire_nl010Ol_o;
			nl01i1i <= wire_nl010ll_o;
			nl01i1l <= wire_nl010lO_o;
			nl01i1O <= wire_nl010Oi_o;
		end
	end
	event nl01i0l_event;
	event nl01i1i_event;
	event nl01i1l_event;
	event nl01i1O_event;
	initial
		#1 ->nl01i0l_event;
	initial
		#1 ->nl01i1i_event;
	initial
		#1 ->nl01i1l_event;
	initial
		#1 ->nl01i1O_event;
	always @(nl01i0l_event)
		nl01i0l <= 1;
	always @(nl01i1i_event)
		nl01i1i <= 1;
	always @(nl01i1l_event)
		nl01i1l <= 1;
	always @(nl01i1O_event)
		nl01i1O <= 1;
	initial
	begin
		nl0i0ll = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nl0i0ll <= 0;
		end
		else if  (n0Oll == 1'b1) 
		begin
			nl0i0ll <= ((((nil10lO & nilOiOl) & (nl1i0OO | nl1i0Oi)) | (~ (nl1i0OO | nl1i0Oi))) & nii00li);
		end
	end
	event nl0i0ll_event;
	initial
		#1 ->nl0i0ll_event;
	always @(nl0i0ll_event)
		nl0i0ll <= 1;
	initial
	begin
		nl0i0Oi = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nl0i0Oi <= 0;
		end
		else if  (wire_nl0i0lO_ENA == 1'b1) 
		begin
			nl0i0Oi <= ((((nil10lO & nilOiOl) & (nl1i0OO | nl1i0Oi)) | (~ (nl1i0OO | nl1i0Oi))) & nii00li);
		end
	end
	assign
		wire_nl0i0lO_ENA = (n0Oll & (~ ni1iili));
	initial
	begin
		nl0i10l = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nl0i10l <= 0;
		end
		else if  (n00il == 1'b1) 
		begin
			nl0i10l <= (nl1i0OO | nl1i0Oi);
		end
	end
	event nl0i10l_event;
	initial
		#1 ->nl0i10l_event;
	always @(nl0i10l_event)
		nl0i10l <= 1;
	initial
	begin
		nl00OlO = 0;
		nl00OOi = 0;
		nl00OOl = 0;
		nl00OOO = 0;
		nl0i11i = 0;
		nl0i11O = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nl00OlO <= 0;
			nl00OOi <= 0;
			nl00OOl <= 0;
			nl00OOO <= 0;
			nl0i11i <= 0;
			nl0i11O <= 0;
		end
		else if  (n01li == 1'b1) 
		begin
			nl00OlO <= nii01li;
			nl00OOi <= nii010i;
			nl00OOl <= nii010l;
			nl00OOO <= nii010O;
			nl0i11i <= nii01ii;
			nl0i11O <= nii01il;
		end
	end
	event nl00OlO_event;
	event nl00OOi_event;
	event nl00OOl_event;
	event nl00OOO_event;
	event nl0i11i_event;
	event nl0i11O_event;
	initial
		#1 ->nl00OlO_event;
	initial
		#1 ->nl00OOi_event;
	initial
		#1 ->nl00OOl_event;
	initial
		#1 ->nl00OOO_event;
	initial
		#1 ->nl0i11i_event;
	initial
		#1 ->nl0i11O_event;
	always @(nl00OlO_event)
		nl00OlO <= 1;
	always @(nl00OOi_event)
		nl00OOi <= 1;
	always @(nl00OOl_event)
		nl00OOl <= 1;
	always @(nl00OOO_event)
		nl00OOO <= 1;
	always @(nl0i11i_event)
		nl0i11i <= 1;
	always @(nl0i11O_event)
		nl0i11O <= 1;
	initial
	begin
		nl0i10O = 0;
		nl0i1ii = 0;
		nl0i1il = 0;
		nl0i1iO = 0;
		nl0i1li = 0;
		nl0i1ll = 0;
		nl0i1lO = 0;
		nl0i1Ol = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nl0i10O <= 0;
			nl0i1ii <= 0;
			nl0i1il <= 0;
			nl0i1iO <= 0;
			nl0i1li <= 0;
			nl0i1ll <= 0;
			nl0i1lO <= 0;
			nl0i1Ol <= 0;
		end
		else if  (ni10O0O == 1'b1) 
		begin
			nl0i10O <= wire_nl0i01i_dataout;
			nl0i1ii <= wire_nl0i01l_dataout;
			nl0i1il <= wire_nl0i01O_dataout;
			nl0i1iO <= wire_nl0i00i_dataout;
			nl0i1li <= wire_nl0i00l_dataout;
			nl0i1ll <= wire_nl0i00O_dataout;
			nl0i1lO <= wire_nl0i0ii_dataout;
			nl0i1Ol <= wire_nl0i1OO_dataout;
		end
	end
	event nl0i10O_event;
	event nl0i1ii_event;
	event nl0i1il_event;
	event nl0i1iO_event;
	event nl0i1li_event;
	event nl0i1ll_event;
	event nl0i1lO_event;
	event nl0i1Ol_event;
	initial
		#1 ->nl0i10O_event;
	initial
		#1 ->nl0i1ii_event;
	initial
		#1 ->nl0i1il_event;
	initial
		#1 ->nl0i1iO_event;
	initial
		#1 ->nl0i1li_event;
	initial
		#1 ->nl0i1ll_event;
	initial
		#1 ->nl0i1lO_event;
	initial
		#1 ->nl0i1Ol_event;
	always @(nl0i10O_event)
		nl0i10O <= 1;
	always @(nl0i1ii_event)
		nl0i1ii <= 1;
	always @(nl0i1il_event)
		nl0i1il <= 1;
	always @(nl0i1iO_event)
		nl0i1iO <= 1;
	always @(nl0i1li_event)
		nl0i1li <= 1;
	always @(nl0i1ll_event)
		nl0i1ll <= 1;
	always @(nl0i1lO_event)
		nl0i1lO <= 1;
	always @(nl0i1Ol_event)
		nl0i1Ol <= 1;
	initial
	begin
		nl0i0OO = 0;
		nl0ii0i = 0;
		nl0ii0l = 0;
		nl0ii0O = 0;
		nl0ii1i = 0;
		nl0ii1l = 0;
		nl0ii1O = 0;
		nl0iiii = 0;
		nl0iiil = 0;
		nl0iili = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nl0i0OO <= 0;
			nl0ii0i <= 0;
			nl0ii0l <= 0;
			nl0ii0O <= 0;
			nl0ii1i <= 0;
			nl0ii1l <= 0;
			nl0ii1O <= 0;
			nl0iiii <= 0;
			nl0iiil <= 0;
			nl0iili <= 0;
		end
		else if  (ni10Oii == 1'b1) 
		begin
			nl0i0OO <= wire_nl0iilO_dataout;
			nl0ii0i <= wire_nl0il1i_dataout;
			nl0ii0l <= wire_nl0il1l_dataout;
			nl0ii0O <= wire_nl0il1O_dataout;
			nl0ii1i <= wire_nl0iiOi_dataout;
			nl0ii1l <= wire_nl0iiOl_dataout;
			nl0ii1O <= wire_nl0iiOO_dataout;
			nl0iiii <= wire_nl0il0i_dataout;
			nl0iiil <= wire_nl0il0l_dataout;
			nl0iili <= wire_nl0iill_dataout;
		end
	end
	event nl0i0OO_event;
	event nl0ii0i_event;
	event nl0ii0l_event;
	event nl0ii0O_event;
	event nl0ii1i_event;
	event nl0ii1l_event;
	event nl0ii1O_event;
	event nl0iiii_event;
	event nl0iiil_event;
	event nl0iili_event;
	initial
		#1 ->nl0i0OO_event;
	initial
		#1 ->nl0ii0i_event;
	initial
		#1 ->nl0ii0l_event;
	initial
		#1 ->nl0ii0O_event;
	initial
		#1 ->nl0ii1i_event;
	initial
		#1 ->nl0ii1l_event;
	initial
		#1 ->nl0ii1O_event;
	initial
		#1 ->nl0iiii_event;
	initial
		#1 ->nl0iiil_event;
	initial
		#1 ->nl0iili_event;
	always @(nl0i0OO_event)
		nl0i0OO <= 1;
	always @(nl0ii0i_event)
		nl0ii0i <= 1;
	always @(nl0ii0l_event)
		nl0ii0l <= 1;
	always @(nl0ii0O_event)
		nl0ii0O <= 1;
	always @(nl0ii1i_event)
		nl0ii1i <= 1;
	always @(nl0ii1l_event)
		nl0ii1l <= 1;
	always @(nl0ii1O_event)
		nl0ii1O <= 1;
	always @(nl0iiii_event)
		nl0iiii <= 1;
	always @(nl0iiil_event)
		nl0iiil <= 1;
	always @(nl0iili_event)
		nl0iili <= 1;
	initial
	begin
		nl0ilil = 0;
		nl0iliO = 0;
		nl0illi = 0;
		nl0illl = 0;
		nl0illO = 0;
		nl0ilOi = 0;
		nl0ilOl = 0;
		nl0ilOO = 0;
		nl0iO1i = 0;
		nl0iO1O = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nl0ilil <= 0;
			nl0iliO <= 0;
			nl0illi <= 0;
			nl0illl <= 0;
			nl0illO <= 0;
			nl0ilOi <= 0;
			nl0ilOl <= 0;
			nl0ilOO <= 0;
			nl0iO1i <= 0;
			nl0iO1O <= 0;
		end
		else if  (ni10Oil == 1'b1) 
		begin
			nl0ilil <= wire_nl0iO0l_dataout;
			nl0iliO <= wire_nl0iO0O_dataout;
			nl0illi <= wire_nl0iOii_dataout;
			nl0illl <= wire_nl0iOil_dataout;
			nl0illO <= wire_nl0iOiO_dataout;
			nl0ilOi <= wire_nl0iOli_dataout;
			nl0ilOl <= wire_nl0iOll_dataout;
			nl0ilOO <= wire_nl0iOlO_dataout;
			nl0iO1i <= wire_nl0iOOi_dataout;
			nl0iO1O <= wire_nl0iO0i_dataout;
		end
	end
	event nl0ilil_event;
	event nl0iliO_event;
	event nl0illi_event;
	event nl0illl_event;
	event nl0illO_event;
	event nl0ilOi_event;
	event nl0ilOl_event;
	event nl0ilOO_event;
	event nl0iO1i_event;
	event nl0iO1O_event;
	initial
		#1 ->nl0ilil_event;
	initial
		#1 ->nl0iliO_event;
	initial
		#1 ->nl0illi_event;
	initial
		#1 ->nl0illl_event;
	initial
		#1 ->nl0illO_event;
	initial
		#1 ->nl0ilOi_event;
	initial
		#1 ->nl0ilOl_event;
	initial
		#1 ->nl0ilOO_event;
	initial
		#1 ->nl0iO1i_event;
	initial
		#1 ->nl0iO1O_event;
	always @(nl0ilil_event)
		nl0ilil <= 1;
	always @(nl0iliO_event)
		nl0iliO <= 1;
	always @(nl0illi_event)
		nl0illi <= 1;
	always @(nl0illl_event)
		nl0illl <= 1;
	always @(nl0illO_event)
		nl0illO <= 1;
	always @(nl0ilOi_event)
		nl0ilOi <= 1;
	always @(nl0ilOl_event)
		nl0ilOl <= 1;
	always @(nl0ilOO_event)
		nl0ilOO <= 1;
	always @(nl0iO1i_event)
		nl0iO1i <= 1;
	always @(nl0iO1O_event)
		nl0iO1O <= 1;
	initial
	begin
		nl0l0il = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nl0l0il <= 0;
		end
		else if  (wire_nl0l0ii_ENA == 1'b1) 
		begin
			nl0l0il <= wire_nl0l00l_o;
		end
	end
	assign
		wire_nl0l0ii_ENA = (n1i1l & (~ ni1iiii));
	event nl0l0il_event;
	initial
		#1 ->nl0l0il_event;
	always @(nl0l0il_event)
		nl0l0il <= 1;
	initial
	begin
		nl0l0Oi = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nl0l0Oi <= 0;
		end
		else if  (wire_nl0l0lO_ENA == 1'b1) 
		begin
			nl0l0Oi <= wire_nl0l0li_o;
		end
	end
	assign
		wire_nl0l0lO_ENA = (n1i1i & (~ ni1iiii));
	event nl0l0Oi_event;
	initial
		#1 ->nl0l0Oi_event;
	always @(nl0l0Oi_event)
		nl0l0Oi <= 1;
	initial
	begin
		nl0li1i = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nl0li1i <= 0;
		end
		else if  (wire_nl0l0OO_ENA == 1'b1) 
		begin
			nl0li1i <= (~ ((((~ nii11OO) & (~ nii11Ol)) & (~ nii11Oi)) & (~ nii11lO)));
		end
	end
	assign
		wire_nl0l0OO_ENA = (n11ii & (~ ni1iiii));
	event nl0li1i_event;
	initial
		#1 ->nl0li1i_event;
	always @(nl0li1i_event)
		nl0li1i <= 1;
	initial
	begin
		nl0l10l = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nl0l10l <= 0;
		end
		else if  (wire_nl0l10i_ENA == 1'b1) 
		begin
			nl0l10l <= (ni10OOl & ni10OOO);
		end
	end
	assign
		wire_nl0l10i_ENA = (n0O1l & (~ ni1iili));
	initial
	begin
		nl0l11l = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nl0l11l <= 0;
		end
		else if  (wire_nl0l11i_ENA == 1'b1) 
		begin
			nl0l11l <= nli1iOO;
		end
	end
	assign
		wire_nl0l11i_ENA = (n0O1l & (~ ni1iili));
	initial
	begin
		nl0l1il = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nl0l1il <= 0;
		end
		else if  (wire_nl0l1ii_ENA == 1'b1) 
		begin
			nl0l1il <= (nl0l10l | nli10iO);
		end
	end
	assign
		wire_nl0l1ii_ENA = (n00ll & (~ ni1iili));
	initial
	begin
		nl0l1ll = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nl0l1ll <= 0;
		end
		else if  (wire_nl0l1li_ENA == 1'b1) 
		begin
			nl0l1ll <= n11ll;
		end
	end
	assign
		wire_nl0l1li_ENA = (n11li & (~ ni1iiii));
	initial
	begin
		nl0l1Oi = 0;
		nl0l1OO = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nl0l1Oi <= 0;
			nl0l1OO <= 0;
		end
		else if  (ni10OiO == 1'b1) 
		begin
			nl0l1Oi <= wire_nl0l01l_dataout;
			nl0l1OO <= wire_nl0l01i_dataout;
		end
	end
	event nl0l1Oi_event;
	event nl0l1OO_event;
	initial
		#1 ->nl0l1Oi_event;
	initial
		#1 ->nl0l1OO_event;
	always @(nl0l1Oi_event)
		nl0l1Oi <= 1;
	always @(nl0l1OO_event)
		nl0l1OO <= 1;
	initial
	begin
		nl0liii = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nl0liii <= 0;
		end
		else if  (wire_nl0li0O_ENA == 1'b1) 
		begin
			nl0liii <= (~ nii1O0i);
		end
	end
	assign
		wire_nl0li0O_ENA = (n110O & (~ ni1iiii));
	event nl0liii_event;
	initial
		#1 ->nl0liii_event;
	always @(nl0liii_event)
		nl0liii <= 1;
	initial
	begin
		nl0li0i = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nl0li0i <= 0;
		end
		else if  (wire_nl0li1O_ENA == 1'b1) 
		begin
			nl0li0i <= ni1i10l;
		end
	end
	assign
		wire_nl0li1O_ENA = (nlOOOO & (~ ni1iiii));
	event nl0li0i_event;
	initial
		#1 ->nl0li0i_event;
	always @(nl0li0i_event)
		nl0li0i <= 1;
	initial
	begin
		nl0lili = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nl0lili <= 0;
		end
		else if  (wire_nl0liiO_ENA == 1'b1) 
		begin
			nl0lili <= nii1iii;
		end
	end
	assign
		wire_nl0liiO_ENA = (n111O & (~ ni1iiii));
	initial
	begin
		nl0lO0i = 0;
		nl0lO0l = 0;
		nl0lO0O = 0;
		nl0lOii = 0;
		nl0lOil = 0;
		nl0lOiO = 0;
		nl0lOli = 0;
		nl0lOll = 0;
		nl0lOlO = 0;
		nl0lOOi = 0;
		nl0lOOO = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nl0lO0i <= 0;
			nl0lO0l <= 0;
			nl0lO0O <= 0;
			nl0lOii <= 0;
			nl0lOil <= 0;
			nl0lOiO <= 0;
			nl0lOli <= 0;
			nl0lOll <= 0;
			nl0lOlO <= 0;
			nl0lOOi <= 0;
			nl0lOOO <= 0;
		end
		else if  (ni10Oli == 1'b1) 
		begin
			nl0lO0i <= wire_nl0O11l_dataout;
			nl0lO0l <= wire_nl0O11O_dataout;
			nl0lO0O <= wire_nl0O10i_dataout;
			nl0lOii <= wire_nl0O10l_dataout;
			nl0lOil <= wire_nl0O10O_dataout;
			nl0lOiO <= wire_nl0O1ii_dataout;
			nl0lOli <= wire_nl0O1il_dataout;
			nl0lOll <= wire_nl0O1iO_dataout;
			nl0lOlO <= wire_nl0O1li_dataout;
			nl0lOOi <= wire_nl0O1ll_dataout;
			nl0lOOO <= wire_nl0O11i_dataout;
		end
	end
	initial
	begin
		nl0O01i = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nl0O01i <= 0;
		end
		else if  (wire_nl0O1OO_ENA == 1'b1) 
		begin
			nl0O01i <= (~ nl0lili);
		end
	end
	assign
		wire_nl0O1OO_ENA = (n110O & (~ ni1iiii));
	initial
	begin
		nl0OiOl = 0;
		nl0OiOO = 0;
		nl0Ol0i = 0;
		nl0Ol0l = 0;
		nl0Ol1i = 0;
		nl0Ol1l = 0;
		nl0Ol1O = 0;
		nl0Olii = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nl0OiOl <= 0;
			nl0OiOO <= 0;
			nl0Ol0i <= 0;
			nl0Ol0l <= 0;
			nl0Ol1i <= 0;
			nl0Ol1l <= 0;
			nl0Ol1O <= 0;
			nl0Olii <= 0;
		end
		else if  (ni1i11i == 1'b1) 
		begin
			nl0OiOl <= wire_nl0Olil_o[2];
			nl0OiOO <= wire_nl0Olil_o[3];
			nl0Ol0i <= wire_nl0Olil_o[7];
			nl0Ol0l <= wire_nl0Olil_o[8];
			nl0Ol1i <= wire_nl0Olil_o[4];
			nl0Ol1l <= wire_nl0Olil_o[5];
			nl0Ol1O <= wire_nl0Olil_o[6];
			nl0Olii <= wire_nl0Olil_o[1];
		end
	end
	event nl0OiOl_event;
	event nl0OiOO_event;
	event nl0Ol0i_event;
	event nl0Ol0l_event;
	event nl0Ol1i_event;
	event nl0Ol1l_event;
	event nl0Ol1O_event;
	event nl0Olii_event;
	initial
		#1 ->nl0OiOl_event;
	initial
		#1 ->nl0OiOO_event;
	initial
		#1 ->nl0Ol0i_event;
	initial
		#1 ->nl0Ol0l_event;
	initial
		#1 ->nl0Ol1i_event;
	initial
		#1 ->nl0Ol1l_event;
	initial
		#1 ->nl0Ol1O_event;
	initial
		#1 ->nl0Olii_event;
	always @(nl0OiOl_event)
		nl0OiOl <= 1;
	always @(nl0OiOO_event)
		nl0OiOO <= 1;
	always @(nl0Ol0i_event)
		nl0Ol0i <= 1;
	always @(nl0Ol0l_event)
		nl0Ol0l <= 1;
	always @(nl0Ol1i_event)
		nl0Ol1i <= 1;
	always @(nl0Ol1l_event)
		nl0Ol1l <= 1;
	always @(nl0Ol1O_event)
		nl0Ol1O <= 1;
	always @(nl0Olii_event)
		nl0Olii <= 1;
	initial
	begin
		nl100iO = 0;
		nl100li = 0;
		nl100ll = 0;
		nl100lO = 0;
		nl100Oi = 0;
		nl100Ol = 0;
		nl100OO = 0;
		nl10i0i = 0;
		nl10i0l = 0;
		nl10i0O = 0;
		nl10i1i = 0;
		nl10i1l = 0;
		nl10i1O = 0;
		nl10iii = 0;
		nl10iil = 0;
		nl10iiO = 0;
		nl10ili = 0;
		nl10ill = 0;
		nl10ilO = 0;
		nl10iOi = 0;
		nl10iOl = 0;
		nl10iOO = 0;
		nl10l1i = 0;
		nl10l1O = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nl100iO <= 0;
			nl100li <= 0;
			nl100ll <= 0;
			nl100lO <= 0;
			nl100Oi <= 0;
			nl100Ol <= 0;
			nl100OO <= 0;
			nl10i0i <= 0;
			nl10i0l <= 0;
			nl10i0O <= 0;
			nl10i1i <= 0;
			nl10i1l <= 0;
			nl10i1O <= 0;
			nl10iii <= 0;
			nl10iil <= 0;
			nl10iiO <= 0;
			nl10ili <= 0;
			nl10ill <= 0;
			nl10ilO <= 0;
			nl10iOi <= 0;
			nl10iOl <= 0;
			nl10iOO <= 0;
			nl10l1i <= 0;
			nl10l1O <= 0;
		end
		else if  (ni101ll == 1'b1) 
		begin
			nl100iO <= wire_nl11Oii_o;
			nl100li <= wire_nl11Oil_o;
			nl100ll <= wire_nl11OiO_o;
			nl100lO <= wire_nl11Oli_o;
			nl100Oi <= wire_nl11Oll_o;
			nl100Ol <= wire_nl11OlO_o;
			nl100OO <= wire_nl11OOi_o;
			nl10i0i <= wire_nl1011l_o;
			nl10i0l <= wire_nl1011O_o;
			nl10i0O <= wire_nl1010i_o;
			nl10i1i <= wire_nl11OOl_o;
			nl10i1l <= wire_nl11OOO_o;
			nl10i1O <= wire_nl1011i_o;
			nl10iii <= wire_nl1010l_o;
			nl10iil <= wire_nl1010O_o;
			nl10iiO <= wire_nl101ii_o;
			nl10ili <= wire_nl101il_o;
			nl10ill <= wire_nl101iO_o;
			nl10ilO <= wire_nl101li_o;
			nl10iOi <= wire_nl101ll_o;
			nl10iOl <= wire_nl101lO_o;
			nl10iOO <= wire_nl101Oi_o;
			nl10l1i <= wire_nl101Ol_o;
			nl10l1O <= wire_nl101OO_o;
		end
	end
	event nl100iO_event;
	event nl100li_event;
	event nl100ll_event;
	event nl100lO_event;
	event nl100Oi_event;
	event nl100Ol_event;
	event nl100OO_event;
	event nl10i0i_event;
	event nl10i0l_event;
	event nl10i0O_event;
	event nl10i1i_event;
	event nl10i1l_event;
	event nl10i1O_event;
	event nl10iii_event;
	event nl10iil_event;
	event nl10iiO_event;
	event nl10ili_event;
	event nl10ill_event;
	event nl10ilO_event;
	event nl10iOi_event;
	event nl10iOl_event;
	event nl10iOO_event;
	event nl10l1i_event;
	event nl10l1O_event;
	initial
		#1 ->nl100iO_event;
	initial
		#1 ->nl100li_event;
	initial
		#1 ->nl100ll_event;
	initial
		#1 ->nl100lO_event;
	initial
		#1 ->nl100Oi_event;
	initial
		#1 ->nl100Ol_event;
	initial
		#1 ->nl100OO_event;
	initial
		#1 ->nl10i0i_event;
	initial
		#1 ->nl10i0l_event;
	initial
		#1 ->nl10i0O_event;
	initial
		#1 ->nl10i1i_event;
	initial
		#1 ->nl10i1l_event;
	initial
		#1 ->nl10i1O_event;
	initial
		#1 ->nl10iii_event;
	initial
		#1 ->nl10iil_event;
	initial
		#1 ->nl10iiO_event;
	initial
		#1 ->nl10ili_event;
	initial
		#1 ->nl10ill_event;
	initial
		#1 ->nl10ilO_event;
	initial
		#1 ->nl10iOi_event;
	initial
		#1 ->nl10iOl_event;
	initial
		#1 ->nl10iOO_event;
	initial
		#1 ->nl10l1i_event;
	initial
		#1 ->nl10l1O_event;
	always @(nl100iO_event)
		nl100iO <= 1;
	always @(nl100li_event)
		nl100li <= 1;
	always @(nl100ll_event)
		nl100ll <= 1;
	always @(nl100lO_event)
		nl100lO <= 1;
	always @(nl100Oi_event)
		nl100Oi <= 1;
	always @(nl100Ol_event)
		nl100Ol <= 1;
	always @(nl100OO_event)
		nl100OO <= 1;
	always @(nl10i0i_event)
		nl10i0i <= 1;
	always @(nl10i0l_event)
		nl10i0l <= 1;
	always @(nl10i0O_event)
		nl10i0O <= 1;
	always @(nl10i1i_event)
		nl10i1i <= 1;
	always @(nl10i1l_event)
		nl10i1l <= 1;
	always @(nl10i1O_event)
		nl10i1O <= 1;
	always @(nl10iii_event)
		nl10iii <= 1;
	always @(nl10iil_event)
		nl10iil <= 1;
	always @(nl10iiO_event)
		nl10iiO <= 1;
	always @(nl10ili_event)
		nl10ili <= 1;
	always @(nl10ill_event)
		nl10ill <= 1;
	always @(nl10ilO_event)
		nl10ilO <= 1;
	always @(nl10iOi_event)
		nl10iOi <= 1;
	always @(nl10iOl_event)
		nl10iOl <= 1;
	always @(nl10iOO_event)
		nl10iOO <= 1;
	always @(nl10l1i_event)
		nl10l1i <= 1;
	always @(nl10l1O_event)
		nl10l1O <= 1;
	initial
	begin
		nl10llO = 0;
		nl10lOO = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nl10llO <= 1;
			nl10lOO <= 1;
		end
		else if  (ni101lO == 1'b1) 
		begin
			nl10llO <= nii1iOO;
			nl10lOO <= nii1l1l;
		end
	end
	event nl10llO_event;
	event nl10lOO_event;
	initial
		#1 ->nl10llO_event;
	initial
		#1 ->nl10lOO_event;
	always @(nl10llO_event)
		nl10llO <= 1;
	always @(nl10lOO_event)
		nl10lOO <= 1;
	initial
	begin
		nl10l0O = 0;
		nl10lii = 0;
		nl10lil = 0;
		nl10liO = 0;
		nl10lli = 0;
		nl10lll = 0;
		nl10lOi = 0;
		nl10O1l = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nl10l0O <= 0;
			nl10lii <= 0;
			nl10lil <= 0;
			nl10liO <= 0;
			nl10lli <= 0;
			nl10lll <= 0;
			nl10lOi <= 0;
			nl10O1l <= 0;
		end
		else if  (ni101lO == 1'b1) 
		begin
			nl10l0O <= nii1iiO;
			nl10lii <= nii1ili;
			nl10lil <= nii1ill;
			nl10liO <= nii1ilO;
			nl10lli <= nii1iOi;
			nl10lll <= nii1iOl;
			nl10lOi <= nii1l1i;
			nl10O1l <= nii1l0i;
		end
	end
	event nl10l0O_event;
	event nl10lii_event;
	event nl10lil_event;
	event nl10liO_event;
	event nl10lli_event;
	event nl10lll_event;
	event nl10lOi_event;
	event nl10O1l_event;
	initial
		#1 ->nl10l0O_event;
	initial
		#1 ->nl10lii_event;
	initial
		#1 ->nl10lil_event;
	initial
		#1 ->nl10liO_event;
	initial
		#1 ->nl10lli_event;
	initial
		#1 ->nl10lll_event;
	initial
		#1 ->nl10lOi_event;
	initial
		#1 ->nl10O1l_event;
	always @(nl10l0O_event)
		nl10l0O <= 1;
	always @(nl10lii_event)
		nl10lii <= 1;
	always @(nl10lil_event)
		nl10lil <= 1;
	always @(nl10liO_event)
		nl10liO <= 1;
	always @(nl10lli_event)
		nl10lli <= 1;
	always @(nl10lll_event)
		nl10lll <= 1;
	always @(nl10lOi_event)
		nl10lOi <= 1;
	always @(nl10O1l_event)
		nl10O1l <= 1;
	initial
	begin
		nl10Oll = 0;
		nl10OOl = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nl10Oll <= 1;
			nl10OOl <= 1;
		end
		else if  (ni101Oi == 1'b1) 
		begin
			nl10Oll <= nii1iOO;
			nl10OOl <= nii1l1l;
		end
	end
	event nl10Oll_event;
	event nl10OOl_event;
	initial
		#1 ->nl10Oll_event;
	initial
		#1 ->nl10OOl_event;
	always @(nl10Oll_event)
		nl10Oll <= 1;
	always @(nl10OOl_event)
		nl10OOl <= 1;
	initial
	begin
		nl10O0l = 0;
		nl10O0O = 0;
		nl10Oii = 0;
		nl10Oil = 0;
		nl10OiO = 0;
		nl10Oli = 0;
		nl10OlO = 0;
		nl1i11i = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nl10O0l <= 0;
			nl10O0O <= 0;
			nl10Oii <= 0;
			nl10Oil <= 0;
			nl10OiO <= 0;
			nl10Oli <= 0;
			nl10OlO <= 0;
			nl1i11i <= 0;
		end
		else if  (ni101Oi == 1'b1) 
		begin
			nl10O0l <= nii1iiO;
			nl10O0O <= nii1ili;
			nl10Oii <= nii1ill;
			nl10Oil <= nii1ilO;
			nl10OiO <= nii1iOi;
			nl10Oli <= nii1iOl;
			nl10OlO <= nii1l1i;
			nl1i11i <= nii1l0i;
		end
	end
	event nl10O0l_event;
	event nl10O0O_event;
	event nl10Oii_event;
	event nl10Oil_event;
	event nl10OiO_event;
	event nl10Oli_event;
	event nl10OlO_event;
	event nl1i11i_event;
	initial
		#1 ->nl10O0l_event;
	initial
		#1 ->nl10O0O_event;
	initial
		#1 ->nl10Oii_event;
	initial
		#1 ->nl10Oil_event;
	initial
		#1 ->nl10OiO_event;
	initial
		#1 ->nl10Oli_event;
	initial
		#1 ->nl10OlO_event;
	initial
		#1 ->nl1i11i_event;
	always @(nl10O0l_event)
		nl10O0l <= 1;
	always @(nl10O0O_event)
		nl10O0O <= 1;
	always @(nl10Oii_event)
		nl10Oii <= 1;
	always @(nl10Oil_event)
		nl10Oil <= 1;
	always @(nl10OiO_event)
		nl10OiO <= 1;
	always @(nl10Oli_event)
		nl10Oli <= 1;
	always @(nl10OlO_event)
		nl10OlO <= 1;
	always @(nl1i11i_event)
		nl1i11i <= 1;
	initial
	begin
		nl1100i = 0;
		nl1100l = 0;
		nl1100O = 0;
		nl1101l = 0;
		nl1101O = 0;
		nl110ii = 0;
		nl110il = 0;
		nl110iO = 0;
		nl110li = 0;
		nl110ll = 0;
		nl110lO = 0;
		nl110Oi = 0;
		nl110Ol = 0;
		nl110OO = 0;
		nl11i0i = 0;
		nl11i0l = 0;
		nl11i0O = 0;
		nl11i1i = 0;
		nl11i1l = 0;
		nl11i1O = 0;
		nl11iii = 0;
		nl11iil = 0;
		nl11iiO = 0;
		nl11ill = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nl1100i <= 0;
			nl1100l <= 0;
			nl1100O <= 0;
			nl1101l <= 0;
			nl1101O <= 0;
			nl110ii <= 0;
			nl110il <= 0;
			nl110iO <= 0;
			nl110li <= 0;
			nl110ll <= 0;
			nl110lO <= 0;
			nl110Oi <= 0;
			nl110Ol <= 0;
			nl110OO <= 0;
			nl11i0i <= 0;
			nl11i0l <= 0;
			nl11i0O <= 0;
			nl11i1i <= 0;
			nl11i1l <= 0;
			nl11i1O <= 0;
			nl11iii <= 0;
			nl11iil <= 0;
			nl11iiO <= 0;
			nl11ill <= 0;
		end
		else if  (ni1010O == 1'b1) 
		begin
			nl1100i <= wire_niOOO1l_o;
			nl1100l <= wire_niOOO1O_o;
			nl1100O <= wire_niOOO0i_o;
			nl1101l <= wire_niOOlOO_o;
			nl1101O <= wire_niOOO1i_o;
			nl110ii <= wire_niOOO0l_o;
			nl110il <= wire_niOOO0O_o;
			nl110iO <= wire_niOOOii_o;
			nl110li <= wire_niOOOil_o;
			nl110ll <= wire_niOOOiO_o;
			nl110lO <= wire_niOOOli_o;
			nl110Oi <= wire_niOOOll_o;
			nl110Ol <= wire_niOOOlO_o;
			nl110OO <= wire_niOOOOi_o;
			nl11i0i <= wire_nl1111l_o;
			nl11i0l <= wire_nl1111O_o;
			nl11i0O <= wire_nl1110i_o;
			nl11i1i <= wire_niOOOOl_o;
			nl11i1l <= wire_niOOOOO_o;
			nl11i1O <= wire_nl1111i_o;
			nl11iii <= wire_nl1110l_o;
			nl11iil <= wire_nl1110O_o;
			nl11iiO <= wire_nl111ii_o;
			nl11ill <= wire_nl111il_o;
		end
	end
	initial
	begin
		nl1i00l = 0;
		nl1i01i = 0;
		nl1i01l = 0;
		nl1i01O = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nl1i00l <= 0;
			nl1i01i <= 0;
			nl1i01l <= 0;
			nl1i01O <= 0;
		end
		else if  (ni101OO == 1'b1) 
		begin
			nl1i00l <= nii1lli;
			nl1i01i <= nii1lii;
			nl1i01l <= nii1lil;
			nl1i01O <= nii1liO;
		end
	end
	event nl1i00l_event;
	event nl1i01i_event;
	event nl1i01l_event;
	event nl1i01O_event;
	initial
		#1 ->nl1i00l_event;
	initial
		#1 ->nl1i01i_event;
	initial
		#1 ->nl1i01l_event;
	initial
		#1 ->nl1i01O_event;
	always @(nl1i00l_event)
		nl1i00l <= 1;
	always @(nl1i01i_event)
		nl1i01i <= 1;
	always @(nl1i01l_event)
		nl1i01l <= 1;
	always @(nl1i01O_event)
		nl1i01O <= 1;
	initial
	begin
		nl1i00O = 0;
		nl1i0ii = 0;
		nl1i0il = 0;
		nl1i0li = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nl1i00O <= 1;
			nl1i0ii <= 1;
			nl1i0il <= 1;
			nl1i0li <= 1;
		end
		else if  (ni101OO == 1'b1) 
		begin
			nl1i00O <= nii1lll;
			nl1i0ii <= nii1llO;
			nl1i0il <= nii1lOi;
			nl1i0li <= nii1lOO;
		end
	end
	event nl1i00O_event;
	event nl1i0ii_event;
	event nl1i0il_event;
	event nl1i0li_event;
	initial
		#1 ->nl1i00O_event;
	initial
		#1 ->nl1i0ii_event;
	initial
		#1 ->nl1i0il_event;
	initial
		#1 ->nl1i0li_event;
	always @(nl1i00O_event)
		nl1i00O <= 1;
	always @(nl1i0ii_event)
		nl1i0ii <= 1;
	always @(nl1i0il_event)
		nl1i0il <= 1;
	always @(nl1i0li_event)
		nl1i0li <= 1;
	initial
	begin
		nl1i0Oi = 0;
		nl1i0OO = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nl1i0Oi <= 0;
			nl1i0OO <= 0;
		end
		else if  (ni1001i == 1'b1) 
		begin
			nl1i0Oi <= wire_niOl0il_q_a[0];
			nl1i0OO <= wire_niOl0il_q_a[1];
		end
	end
	event nl1i0Oi_event;
	event nl1i0OO_event;
	initial
		#1 ->nl1i0Oi_event;
	initial
		#1 ->nl1i0OO_event;
	always @(nl1i0Oi_event)
		nl1i0Oi <= 1;
	always @(nl1i0OO_event)
		nl1i0OO <= 1;
	initial
	begin
		nl1i10i = 0;
		nl1i10l = 0;
		nl1i10O = 0;
		nl1i1il = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nl1i10i <= 0;
			nl1i10l <= 0;
			nl1i10O <= 0;
			nl1i1il <= 0;
		end
		else if  (ni101Ol == 1'b1) 
		begin
			nl1i10i <= nii1lii;
			nl1i10l <= nii1lil;
			nl1i10O <= nii1liO;
			nl1i1il <= nii1lli;
		end
	end
	event nl1i10i_event;
	event nl1i10l_event;
	event nl1i10O_event;
	event nl1i1il_event;
	initial
		#1 ->nl1i10i_event;
	initial
		#1 ->nl1i10l_event;
	initial
		#1 ->nl1i10O_event;
	initial
		#1 ->nl1i1il_event;
	always @(nl1i10i_event)
		nl1i10i <= 1;
	always @(nl1i10l_event)
		nl1i10l <= 1;
	always @(nl1i10O_event)
		nl1i10O <= 1;
	always @(nl1i1il_event)
		nl1i1il <= 1;
	initial
	begin
		nl1i1iO = 0;
		nl1i1li = 0;
		nl1i1ll = 0;
		nl1i1Oi = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nl1i1iO <= 1;
			nl1i1li <= 1;
			nl1i1ll <= 1;
			nl1i1Oi <= 1;
		end
		else if  (ni101Ol == 1'b1) 
		begin
			nl1i1iO <= nii1lll;
			nl1i1li <= nii1llO;
			nl1i1ll <= nii1lOi;
			nl1i1Oi <= nii1lOO;
		end
	end
	event nl1i1iO_event;
	event nl1i1li_event;
	event nl1i1ll_event;
	event nl1i1Oi_event;
	initial
		#1 ->nl1i1iO_event;
	initial
		#1 ->nl1i1li_event;
	initial
		#1 ->nl1i1ll_event;
	initial
		#1 ->nl1i1Oi_event;
	always @(nl1i1iO_event)
		nl1i1iO <= 1;
	always @(nl1i1li_event)
		nl1i1li <= 1;
	always @(nl1i1ll_event)
		nl1i1ll <= 1;
	always @(nl1i1Oi_event)
		nl1i1Oi <= 1;
	initial
	begin
		nl1ii0i = 0;
		nl1ii0l = 0;
		nl1ii0O = 0;
		nl1ii1l = 0;
		nl1ii1O = 0;
		nl1iiii = 0;
		nl1iiil = 0;
		nl1iili = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nl1ii0i <= 0;
			nl1ii0l <= 0;
			nl1ii0O <= 0;
			nl1ii1l <= 0;
			nl1ii1O <= 0;
			nl1iiii <= 0;
			nl1iiil <= 0;
			nl1iili <= 0;
		end
		else if  (ni1001l == 1'b1) 
		begin
			nl1ii0i <= nl1100l;
			nl1ii0l <= nl1100O;
			nl1ii0O <= nl110ii;
			nl1ii1l <= nl1101O;
			nl1ii1O <= nl1100i;
			nl1iiii <= nl110il;
			nl1iiil <= nl110iO;
			nl1iili <= nl1101l;
		end
	end
	initial
	begin
		nl1iilO = 0;
		nl1iiOi = 0;
		nl1iiOl = 0;
		nl1iiOO = 0;
		nl1il0l = 0;
		nl1il1i = 0;
		nl1il1l = 0;
		nl1il1O = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nl1iilO <= 0;
			nl1iiOi <= 0;
			nl1iiOl <= 0;
			nl1iiOO <= 0;
			nl1il0l <= 0;
			nl1il1i <= 0;
			nl1il1l <= 0;
			nl1il1O <= 0;
		end
		else if  (ni1001O == 1'b1) 
		begin
			nl1iilO <= nl110ll;
			nl1iiOi <= nl110lO;
			nl1iiOl <= nl110Oi;
			nl1iiOO <= nl110Ol;
			nl1il0l <= nl110li;
			nl1il1i <= nl110OO;
			nl1il1l <= nl11i1i;
			nl1il1O <= nl11i1l;
		end
	end
	initial
	begin
		nl1ilii = 0;
		nl1ilil = 0;
		nl1iliO = 0;
		nl1illi = 0;
		nl1illl = 0;
		nl1illO = 0;
		nl1ilOi = 0;
		nl1ilOO = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nl1ilii <= 0;
			nl1ilil <= 0;
			nl1iliO <= 0;
			nl1illi <= 0;
			nl1illl <= 0;
			nl1illO <= 0;
			nl1ilOi <= 0;
			nl1ilOO <= 0;
		end
		else if  (ni1000i == 1'b1) 
		begin
			nl1ilii <= nl11i0i;
			nl1ilil <= nl11i0l;
			nl1iliO <= nl11i0O;
			nl1illi <= nl11iii;
			nl1illl <= nl11iil;
			nl1illO <= nl11iiO;
			nl1ilOi <= nl11ill;
			nl1ilOO <= nl11i1O;
		end
	end
	event nl1ilii_event;
	event nl1ilil_event;
	event nl1iliO_event;
	event nl1illi_event;
	event nl1illl_event;
	event nl1illO_event;
	event nl1ilOi_event;
	event nl1ilOO_event;
	initial
		#1 ->nl1ilii_event;
	initial
		#1 ->nl1ilil_event;
	initial
		#1 ->nl1iliO_event;
	initial
		#1 ->nl1illi_event;
	initial
		#1 ->nl1illl_event;
	initial
		#1 ->nl1illO_event;
	initial
		#1 ->nl1ilOi_event;
	initial
		#1 ->nl1ilOO_event;
	always @(nl1ilii_event)
		nl1ilii <= 1;
	always @(nl1ilil_event)
		nl1ilil <= 1;
	always @(nl1iliO_event)
		nl1iliO <= 1;
	always @(nl1illi_event)
		nl1illi <= 1;
	always @(nl1illl_event)
		nl1illl <= 1;
	always @(nl1illO_event)
		nl1illO <= 1;
	always @(nl1ilOi_event)
		nl1ilOi <= 1;
	always @(nl1ilOO_event)
		nl1ilOO <= 1;
	initial
	begin
		nl1iO0i = 0;
		nl1iO0l = 0;
		nl1iO0O = 0;
		nl1iO1l = 0;
		nl1iO1O = 0;
		nl1iOii = 0;
		nl1iOil = 0;
		nl1iOli = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nl1iO0i <= 0;
			nl1iO0l <= 0;
			nl1iO0O <= 0;
			nl1iO1l <= 0;
			nl1iO1O <= 0;
			nl1iOii <= 0;
			nl1iOil <= 0;
			nl1iOli <= 0;
		end
		else if  (ni1000l == 1'b1) 
		begin
			nl1iO0i <= wire_nl1iOll_o[11];
			nl1iO0l <= wire_nl1iOll_o[12];
			nl1iO0O <= wire_nl1iOll_o[13];
			nl1iO1l <= wire_nl1iOll_o[9];
			nl1iO1O <= wire_nl1iOll_o[10];
			nl1iOii <= wire_nl1iOll_o[14];
			nl1iOil <= wire_nl1iOll_o[15];
			nl1iOli <= wire_nl1iOll_o[16];
		end
	end
	event nl1iO0i_event;
	event nl1iO0l_event;
	event nl1iO0O_event;
	event nl1iO1l_event;
	event nl1iO1O_event;
	event nl1iOii_event;
	event nl1iOil_event;
	event nl1iOli_event;
	initial
		#1 ->nl1iO0i_event;
	initial
		#1 ->nl1iO0l_event;
	initial
		#1 ->nl1iO0O_event;
	initial
		#1 ->nl1iO1l_event;
	initial
		#1 ->nl1iO1O_event;
	initial
		#1 ->nl1iOii_event;
	initial
		#1 ->nl1iOil_event;
	initial
		#1 ->nl1iOli_event;
	always @(nl1iO0i_event)
		nl1iO0i <= 1;
	always @(nl1iO0l_event)
		nl1iO0l <= 1;
	always @(nl1iO0O_event)
		nl1iO0O <= 1;
	always @(nl1iO1l_event)
		nl1iO1l <= 1;
	always @(nl1iO1O_event)
		nl1iO1O <= 1;
	always @(nl1iOii_event)
		nl1iOii <= 1;
	always @(nl1iOil_event)
		nl1iOil <= 1;
	always @(nl1iOli_event)
		nl1iOli <= 1;
	initial
	begin
		nl1l01l = 0;
		nl1l1iO = 0;
		nl1l1li = 0;
		nl1l1ll = 0;
		nl1l1lO = 0;
		nl1l1Oi = 0;
		nl1l1Ol = 0;
		nl1l1OO = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nl1l01l <= 0;
			nl1l1iO <= 0;
			nl1l1li <= 0;
			nl1l1ll <= 0;
			nl1l1lO <= 0;
			nl1l1Oi <= 0;
			nl1l1Ol <= 0;
			nl1l1OO <= 0;
		end
		else if  (ni100ii == 1'b1) 
		begin
			nl1l01l <= wire_nl1l01O_o[16];
			nl1l1iO <= wire_nl1l01O_o[9];
			nl1l1li <= wire_nl1l01O_o[10];
			nl1l1ll <= wire_nl1l01O_o[11];
			nl1l1lO <= wire_nl1l01O_o[12];
			nl1l1Oi <= wire_nl1l01O_o[13];
			nl1l1Ol <= wire_nl1l01O_o[14];
			nl1l1OO <= wire_nl1l01O_o[15];
		end
	end
	event nl1l01l_event;
	event nl1l1iO_event;
	event nl1l1li_event;
	event nl1l1ll_event;
	event nl1l1lO_event;
	event nl1l1Oi_event;
	event nl1l1Ol_event;
	event nl1l1OO_event;
	initial
		#1 ->nl1l01l_event;
	initial
		#1 ->nl1l1iO_event;
	initial
		#1 ->nl1l1li_event;
	initial
		#1 ->nl1l1ll_event;
	initial
		#1 ->nl1l1lO_event;
	initial
		#1 ->nl1l1Oi_event;
	initial
		#1 ->nl1l1Ol_event;
	initial
		#1 ->nl1l1OO_event;
	always @(nl1l01l_event)
		nl1l01l <= 1;
	always @(nl1l1iO_event)
		nl1l1iO <= 1;
	always @(nl1l1li_event)
		nl1l1li <= 1;
	always @(nl1l1ll_event)
		nl1l1ll <= 1;
	always @(nl1l1lO_event)
		nl1l1lO <= 1;
	always @(nl1l1Oi_event)
		nl1l1Oi <= 1;
	always @(nl1l1Ol_event)
		nl1l1Ol <= 1;
	always @(nl1l1OO_event)
		nl1l1OO <= 1;
	initial
	begin
		nl1iOOi = 0;
		nl1iOOl = 0;
		nl1iOOO = 0;
		nl1l10i = 0;
		nl1l10O = 0;
		nl1l11i = 0;
		nl1l11l = 0;
		nl1l11O = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nl1iOOi <= 0;
			nl1iOOl <= 0;
			nl1iOOO <= 0;
			nl1l10i <= 0;
			nl1l10O <= 0;
			nl1l11i <= 0;
			nl1l11l <= 0;
			nl1l11O <= 0;
		end
		else if  (ni1000O == 1'b1) 
		begin
			nl1iOOi <= wire_nl1l1ii_o[9];
			nl1iOOl <= wire_nl1l1ii_o[10];
			nl1iOOO <= wire_nl1l1ii_o[11];
			nl1l10i <= wire_nl1l1ii_o[15];
			nl1l10O <= wire_nl1l1ii_o[16];
			nl1l11i <= wire_nl1l1ii_o[12];
			nl1l11l <= wire_nl1l1ii_o[13];
			nl1l11O <= wire_nl1l1ii_o[14];
		end
	end
	event nl1iOOi_event;
	event nl1iOOl_event;
	event nl1iOOO_event;
	event nl1l10i_event;
	event nl1l10O_event;
	event nl1l11i_event;
	event nl1l11l_event;
	event nl1l11O_event;
	initial
		#1 ->nl1iOOi_event;
	initial
		#1 ->nl1iOOl_event;
	initial
		#1 ->nl1iOOO_event;
	initial
		#1 ->nl1l10i_event;
	initial
		#1 ->nl1l10O_event;
	initial
		#1 ->nl1l11i_event;
	initial
		#1 ->nl1l11l_event;
	initial
		#1 ->nl1l11O_event;
	always @(nl1iOOi_event)
		nl1iOOi <= 1;
	always @(nl1iOOl_event)
		nl1iOOl <= 1;
	always @(nl1iOOO_event)
		nl1iOOO <= 1;
	always @(nl1l10i_event)
		nl1l10i <= 1;
	always @(nl1l10O_event)
		nl1l10O <= 1;
	always @(nl1l11i_event)
		nl1l11i <= 1;
	always @(nl1l11l_event)
		nl1l11l <= 1;
	always @(nl1l11O_event)
		nl1l11O <= 1;
	initial
	begin
		nl1llll = 0;
		nl1lllO = 0;
		nl1llOi = 0;
		nl1llOl = 0;
		nl1llOO = 0;
		nl1lO0i = 0;
		nl1lO1i = 0;
		nl1lO1l = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nl1llll <= 0;
			nl1lllO <= 0;
			nl1llOi <= 0;
			nl1llOl <= 0;
			nl1llOO <= 0;
			nl1lO0i <= 0;
			nl1lO1i <= 0;
			nl1lO1l <= 0;
		end
		else if  (ni100il == 1'b1) 
		begin
			nl1llll <= wire_nl1lO0O_dataout;
			nl1lllO <= wire_nl1lOii_dataout;
			nl1llOi <= wire_nl1lOil_dataout;
			nl1llOl <= wire_nl1lOiO_dataout;
			nl1llOO <= wire_nl1lOli_dataout;
			nl1lO0i <= wire_nl1lO0l_dataout;
			nl1lO1i <= wire_nl1lOll_dataout;
			nl1lO1l <= wire_nl1lOlO_dataout;
		end
	end
	initial
	begin
		nl1O00i = 0;
		nl1O00O = 0;
		nl1O01i = 0;
		nl1O01l = 0;
		nl1O01O = 0;
		nl1O1lO = 0;
		nl1O1Oi = 0;
		nl1O1Ol = 0;
		nl1O1OO = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nl1O00i <= 0;
			nl1O00O <= 0;
			nl1O01i <= 0;
			nl1O01l <= 0;
			nl1O01O <= 0;
			nl1O1lO <= 0;
			nl1O1Oi <= 0;
			nl1O1Ol <= 0;
			nl1O1OO <= 0;
		end
		else if  (ni100li == 1'b1) 
		begin
			nl1O00i <= wire_nl1O0OO_dataout;
			nl1O00O <= wire_nl1O0ii_dataout;
			nl1O01i <= wire_nl1O0lO_dataout;
			nl1O01l <= wire_nl1O0Oi_dataout;
			nl1O01O <= wire_nl1O0Ol_dataout;
			nl1O1lO <= wire_nl1O0il_dataout;
			nl1O1Oi <= wire_nl1O0iO_dataout;
			nl1O1Ol <= wire_nl1O0li_dataout;
			nl1O1OO <= wire_nl1O0ll_dataout;
		end
	end
	event nl1O00i_event;
	event nl1O00O_event;
	event nl1O01i_event;
	event nl1O01l_event;
	event nl1O01O_event;
	event nl1O1lO_event;
	event nl1O1Oi_event;
	event nl1O1Ol_event;
	event nl1O1OO_event;
	initial
		#1 ->nl1O00i_event;
	initial
		#1 ->nl1O00O_event;
	initial
		#1 ->nl1O01i_event;
	initial
		#1 ->nl1O01l_event;
	initial
		#1 ->nl1O01O_event;
	initial
		#1 ->nl1O1lO_event;
	initial
		#1 ->nl1O1Oi_event;
	initial
		#1 ->nl1O1Ol_event;
	initial
		#1 ->nl1O1OO_event;
	always @(nl1O00i_event)
		nl1O00i <= 1;
	always @(nl1O00O_event)
		nl1O00O <= 1;
	always @(nl1O01i_event)
		nl1O01i <= 1;
	always @(nl1O01l_event)
		nl1O01l <= 1;
	always @(nl1O01O_event)
		nl1O01O <= 1;
	always @(nl1O1lO_event)
		nl1O1lO <= 1;
	always @(nl1O1Oi_event)
		nl1O1Oi <= 1;
	always @(nl1O1Ol_event)
		nl1O1Ol <= 1;
	always @(nl1O1OO_event)
		nl1O1OO <= 1;
	initial
	begin
		nl1O10i = 0;
		nl1O10l = 0;
		nl1O10O = 0;
		nl1O11i = 0;
		nl1O11l = 0;
		nl1O11O = 0;
		nl1O1ii = 0;
		nl1O1il = 0;
		nl1O1li = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nl1O10i <= 0;
			nl1O10l <= 0;
			nl1O10O <= 0;
			nl1O11i <= 0;
			nl1O11l <= 0;
			nl1O11O <= 0;
			nl1O1ii <= 0;
			nl1O1il <= 0;
			nl1O1li <= 0;
		end
		else if  (ni100iO == 1'b1) 
		begin
			nl1O10i <= (nl1llOi & (~ ni1i10i));
			nl1O10l <= (nl1llOl & (~ ni1i10i));
			nl1O10O <= (nl1llOO & (~ ni1i10i));
			nl1O11i <= (nl1lO0i & (~ ni1i10i));
			nl1O11l <= (nl1llll & (~ ni1i10i));
			nl1O11O <= (nl1lllO & (~ ni1i10i));
			nl1O1ii <= (nl1lO1i & (~ ni1i10i));
			nl1O1il <= (nl1lO1l & (~ ni1i10i));
			nl1O1li <= ni1i10i;
		end
	end
	event nl1O10i_event;
	event nl1O10l_event;
	event nl1O10O_event;
	event nl1O11i_event;
	event nl1O11l_event;
	event nl1O11O_event;
	event nl1O1ii_event;
	event nl1O1il_event;
	event nl1O1li_event;
	initial
		#1 ->nl1O10i_event;
	initial
		#1 ->nl1O10l_event;
	initial
		#1 ->nl1O10O_event;
	initial
		#1 ->nl1O11i_event;
	initial
		#1 ->nl1O11l_event;
	initial
		#1 ->nl1O11O_event;
	initial
		#1 ->nl1O1ii_event;
	initial
		#1 ->nl1O1il_event;
	initial
		#1 ->nl1O1li_event;
	always @(nl1O10i_event)
		nl1O10i <= 1;
	always @(nl1O10l_event)
		nl1O10l <= 1;
	always @(nl1O10O_event)
		nl1O10O <= 1;
	always @(nl1O11i_event)
		nl1O11i <= 1;
	always @(nl1O11l_event)
		nl1O11l <= 1;
	always @(nl1O11O_event)
		nl1O11O <= 1;
	always @(nl1O1ii_event)
		nl1O1ii <= 1;
	always @(nl1O1il_event)
		nl1O1il <= 1;
	always @(nl1O1li_event)
		nl1O1li <= 1;
	initial
	begin
		niiilOO = 0;
		nil0O1l = 0;
		niO11OO = 0;
		nl1Oi0i = 0;
		nl1Oiil = 0;
		nl1Oili = 0;
		nl1OiOl = 0;
		nl1Ol0l = 0;
		nl1Ol1i = 0;
		nl1Olii = 0;
		nl1Olll = 0;
		nl1OlOi = 0;
		nl1OO0i = 0;
		nl1OO1l = 0;
		nl1OOiO = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			niiilOO <= 0;
			nil0O1l <= 0;
			niO11OO <= 0;
			nl1Oi0i <= 0;
			nl1Oiil <= 0;
			nl1Oili <= 0;
			nl1OiOl <= 0;
			nl1Ol0l <= 0;
			nl1Ol1i <= 0;
			nl1Olii <= 0;
			nl1Olll <= 0;
			nl1OlOi <= 0;
			nl1OO0i <= 0;
			nl1OO1l <= 0;
			nl1OOiO <= 0;
		end
		else if  (ni1iili == 1'b0) 
		begin
			niiilOO <= ni1il1i;
			nil0O1l <= ni1il1i;
			niO11OO <= ni1il1i;
			nl1Oi0i <= nl1Oiil;
			nl1Oiil <= n010l;
			nl1Oili <= nl1OiOl;
			nl1OiOl <= n010l;
			nl1Ol0l <= n010l;
			nl1Ol1i <= nl1Ol0l;
			nl1Olii <= nl1Olll;
			nl1Olll <= n010l;
			nl1OlOi <= nl1OO1l;
			nl1OO0i <= nl1OOiO;
			nl1OO1l <= n010l;
			nl1OOiO <= n010l;
		end
	end
	initial
	begin
		nl1OOll = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nl1OOll <= 0;
		end
		else if  (wire_nl1OOli_ENA == 1'b1) 
		begin
			nl1OOll <= (((((~ (wire_nl0OOii_o[11] | ni1i11l)) & (wire_nli110l_o[11] | ni1i11O)) & (~ wire_nli110O_o[9])) & wire_nli11ii_o[9]) & (nl1i0OO | nl1i0Oi));
		end
	end
	assign
		wire_nl1OOli_ENA = (n0O1l & (~ ni1iili));
	initial
	begin
		nl1OOOl = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nl1OOOl <= 0;
		end
		else if  (wire_nl1OOOi_ENA == 1'b1) 
		begin
			nl1OOOl <= ni1il1i;
		end
	end
	assign
		wire_nl1OOOi_ENA = (n0O1l & (~ ni1iili));
	initial
	begin
		nli000l = 0;
		nli001i = 0;
		nli001l = 0;
		nli001O = 0;
		nli01lO = 0;
		nli01Oi = 0;
		nli01Ol = 0;
		nli01OO = 0;
	end
	always @ ( posedge clock or  negedge wire_nli000i_CLRN)
	begin
		if (wire_nli000i_CLRN == 1'b0) 
		begin
			nli000l <= 0;
			nli001i <= 0;
			nli001l <= 0;
			nli001O <= 0;
			nli01lO <= 0;
			nli01Oi <= 0;
			nli01Ol <= 0;
			nli01OO <= 0;
		end
		else if  (ni1i00i == 1'b1) 
		begin
			nli000l <= nl10iiO;
			nli001i <= nl10i0O;
			nli001l <= nl10iii;
			nli001O <= nl10iil;
			nli01lO <= nl10i1l;
			nli01Oi <= nl10i1O;
			nli01Ol <= nl10i0i;
			nli01OO <= nl10i0l;
		end
	end
	assign
		wire_nli000i_CLRN = ((ni1i01O66 ^ ni1i01O65) & (~ reset));
	event nli000l_event;
	event nli001i_event;
	event nli001l_event;
	event nli001O_event;
	event nli01lO_event;
	event nli01Oi_event;
	event nli01Ol_event;
	event nli01OO_event;
	initial
		#1 ->nli000l_event;
	initial
		#1 ->nli001i_event;
	initial
		#1 ->nli001l_event;
	initial
		#1 ->nli001O_event;
	initial
		#1 ->nli01lO_event;
	initial
		#1 ->nli01Oi_event;
	initial
		#1 ->nli01Ol_event;
	initial
		#1 ->nli01OO_event;
	always @(nli000l_event)
		nli000l <= 1;
	always @(nli001i_event)
		nli001i <= 1;
	always @(nli001l_event)
		nli001l <= 1;
	always @(nli001O_event)
		nli001O <= 1;
	always @(nli01lO_event)
		nli01lO <= 1;
	always @(nli01Oi_event)
		nli01Oi <= 1;
	always @(nli01Ol_event)
		nli01Ol <= 1;
	always @(nli01OO_event)
		nli01OO <= 1;
	initial
	begin
		nli00ii = 0;
		nli00il = 0;
		nli00iO = 0;
		nli00li = 0;
		nli00ll = 0;
		nli00lO = 0;
		nli00Oi = 0;
		nli00OO = 0;
	end
	always @ (clock or wire_nli00Ol_PRN or wire_nli00Ol_CLRN)
	begin
		if (wire_nli00Ol_PRN == 1'b0) 
		begin
			nli00ii <= 1;
			nli00il <= 1;
			nli00iO <= 1;
			nli00li <= 1;
			nli00ll <= 1;
			nli00lO <= 1;
			nli00Oi <= 1;
			nli00OO <= 1;
		end
		else if  (wire_nli00Ol_CLRN == 1'b0) 
		begin
			nli00ii <= 0;
			nli00il <= 0;
			nli00iO <= 0;
			nli00li <= 0;
			nli00ll <= 0;
			nli00lO <= 0;
			nli00Oi <= 0;
			nli00OO <= 0;
		end
		else if  (ni1i0ii == 1'b1) 
		if (clock != nli00Ol_clk_prev && clock == 1'b1) 
		begin
			nli00ii <= nl100iO;
			nli00il <= nl100li;
			nli00iO <= nl100ll;
			nli00li <= nl100lO;
			nli00ll <= nl100Oi;
			nli00lO <= nl100Ol;
			nli00Oi <= nl100OO;
			nli00OO <= nl10i1i;
		end
		nli00Ol_clk_prev <= clock;
	end
	assign
		wire_nli00Ol_CLRN = ((ni1i00O62 ^ ni1i00O61) & (~ reset)),
		wire_nli00Ol_PRN = (ni1i00l64 ^ ni1i00l63);
	initial
	begin
		nli010i = 0;
		nli010l = 0;
		nli010O = 0;
		nli011l = 0;
		nli011O = 0;
		nli01ii = 0;
		nli01il = 0;
		nli01li = 0;
	end
	always @ (clock or wire_nli01iO_PRN or reset)
	begin
		if (wire_nli01iO_PRN == 1'b0) 
		begin
			nli010i <= 1;
			nli010l <= 1;
			nli010O <= 1;
			nli011l <= 1;
			nli011O <= 1;
			nli01ii <= 1;
			nli01il <= 1;
			nli01li <= 1;
		end
		else if  (reset == 1'b1) 
		begin
			nli010i <= 0;
			nli010l <= 0;
			nli010O <= 0;
			nli011l <= 0;
			nli011O <= 0;
			nli01ii <= 0;
			nli01il <= 0;
			nli01li <= 0;
		end
		else if  (ni1i01l == 1'b1) 
		if (clock != nli01iO_clk_prev && clock == 1'b1) 
		begin
			nli010i <= nl10ilO;
			nli010l <= nl10iOi;
			nli010O <= nl10iOl;
			nli011l <= nl10ili;
			nli011O <= nl10ill;
			nli01ii <= nl10iOO;
			nli01il <= nl10l1i;
			nli01li <= nl10l1O;
		end
		nli01iO_clk_prev <= clock;
	end
	assign
		wire_nli01iO_PRN = (ni1i01i68 ^ ni1i01i67);
	initial
	begin
		nli0i0i = 0;
		nli0i0l = 0;
		nli0i0O = 0;
		nli0i1l = 0;
		nli0i1O = 0;
		nli0iii = 0;
		nli0iil = 0;
		nli0ili = 0;
	end
	always @ (clock or wire_nli0iiO_PRN or wire_nli0iiO_CLRN)
	begin
		if (wire_nli0iiO_PRN == 1'b0) 
		begin
			nli0i0i <= 1;
			nli0i0l <= 1;
			nli0i0O <= 1;
			nli0i1l <= 1;
			nli0i1O <= 1;
			nli0iii <= 1;
			nli0iil <= 1;
			nli0ili <= 1;
		end
		else if  (wire_nli0iiO_CLRN == 1'b0) 
		begin
			nli0i0i <= 0;
			nli0i0l <= 0;
			nli0i0O <= 0;
			nli0i1l <= 0;
			nli0i1O <= 0;
			nli0iii <= 0;
			nli0iil <= 0;
			nli0ili <= 0;
		end
		else if  (ni1i0li == 1'b1) 
		if (clock != nli0iiO_clk_prev && clock == 1'b1) 
		begin
			nli0i0i <= nli1OiO;
			nli0i0l <= nli1Oli;
			nli0i0O <= nli1Oll;
			nli0i1l <= nli1Oii;
			nli0i1O <= nli1Oil;
			nli0iii <= nli1OlO;
			nli0iil <= nli1OOi;
			nli0ili <= nli1OOO;
		end
		nli0iiO_clk_prev <= clock;
	end
	assign
		wire_nli0iiO_CLRN = ((ni1i0iO58 ^ ni1i0iO57) & (~ reset)),
		wire_nli0iiO_PRN = (ni1i0il60 ^ ni1i0il59);
	event nli0i0i_event;
	event nli0i0l_event;
	event nli0i0O_event;
	event nli0i1l_event;
	event nli0i1O_event;
	event nli0iii_event;
	event nli0iil_event;
	event nli0ili_event;
	initial
		#1 ->nli0i0i_event;
	initial
		#1 ->nli0i0l_event;
	initial
		#1 ->nli0i0O_event;
	initial
		#1 ->nli0i1l_event;
	initial
		#1 ->nli0i1O_event;
	initial
		#1 ->nli0iii_event;
	initial
		#1 ->nli0iil_event;
	initial
		#1 ->nli0ili_event;
	always @(nli0i0i_event)
		nli0i0i <= 1;
	always @(nli0i0l_event)
		nli0i0l <= 1;
	always @(nli0i0O_event)
		nli0i0O <= 1;
	always @(nli0i1l_event)
		nli0i1l <= 1;
	always @(nli0i1O_event)
		nli0i1O <= 1;
	always @(nli0iii_event)
		nli0iii <= 1;
	always @(nli0iil_event)
		nli0iil <= 1;
	always @(nli0ili_event)
		nli0ili <= 1;
	initial
	begin
		nli0ilO = 0;
		nli0iOi = 0;
		nli0iOl = 0;
		nli0iOO = 0;
		nli0l0l = 0;
		nli0l1i = 0;
		nli0l1l = 0;
		nli0l1O = 0;
	end
	always @ ( posedge clock or  negedge wire_nli0l0i_CLRN)
	begin
		if (wire_nli0l0i_CLRN == 1'b0) 
		begin
			nli0ilO <= 0;
			nli0iOi <= 0;
			nli0iOl <= 0;
			nli0iOO <= 0;
			nli0l0l <= 0;
			nli0l1i <= 0;
			nli0l1l <= 0;
			nli0l1O <= 0;
		end
		else if  (ni1i0lO == 1'b1) 
		begin
			nli0ilO <= nli1l1l;
			nli0iOi <= nli1l1O;
			nli0iOl <= nli1l0i;
			nli0iOO <= nli1l0l;
			nli0l0l <= nli1lli;
			nli0l1i <= nli1l0O;
			nli0l1l <= nli1lii;
			nli0l1O <= nli1lil;
		end
	end
	assign
		wire_nli0l0i_CLRN = ((ni1i0ll56 ^ ni1i0ll55) & (~ reset));
	initial
	begin
		nli0lii = 0;
		nli0lil = 0;
		nli0liO = 0;
		nli0lli = 0;
		nli0lll = 0;
		nli0llO = 0;
		nli0lOi = 0;
		nli0lOO = 0;
	end
	always @ (clock or wire_nli0lOl_PRN or wire_nli0lOl_CLRN)
	begin
		if (wire_nli0lOl_PRN == 1'b0) 
		begin
			nli0lii <= 1;
			nli0lil <= 1;
			nli0liO <= 1;
			nli0lli <= 1;
			nli0lll <= 1;
			nli0llO <= 1;
			nli0lOi <= 1;
			nli0lOO <= 1;
		end
		else if  (wire_nli0lOl_CLRN == 1'b0) 
		begin
			nli0lii <= 0;
			nli0lil <= 0;
			nli0liO <= 0;
			nli0lli <= 0;
			nli0lll <= 0;
			nli0llO <= 0;
			nli0lOi <= 0;
			nli0lOO <= 0;
		end
		else if  (ni1i0OO == 1'b1) 
		if (clock != nli0lOl_clk_prev && clock == 1'b1) 
		begin
			nli0lii <= nli1llO;
			nli0lil <= nli1lOi;
			nli0liO <= nli1lOl;
			nli0lli <= nli1lOO;
			nli0lll <= nli1O1i;
			nli0llO <= nli1O1l;
			nli0lOi <= nli1O1O;
			nli0lOO <= nli1O0l;
		end
		nli0lOl_clk_prev <= clock;
	end
	assign
		wire_nli0lOl_CLRN = ((ni1i0Ol52 ^ ni1i0Ol51) & (~ reset)),
		wire_nli0lOl_PRN = (ni1i0Oi54 ^ ni1i0Oi53);
	initial
	begin
		nli100O = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nli100O <= 0;
		end
		else if  (wire_nli100l_ENA == 1'b1) 
		begin
			nli100O <= nl1OOll;
		end
	end
	assign
		wire_nli100l_ENA = (n00ll & (~ ni1iili));
	initial
	begin
		nli101O = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nli101O <= 0;
		end
		else if  (wire_nli101l_ENA == 1'b1) 
		begin
			nli101O <= nl0l11l;
		end
	end
	assign
		wire_nli101l_ENA = (n00ll & (~ ni1iili));
	event nli101O_event;
	initial
		#1 ->nli101O_event;
	always @(nli101O_event)
		nli101O <= 1;
	initial
	begin
		nli10iO = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nli10iO <= 0;
		end
		else if  (wire_nli10il_ENA == 1'b1) 
		begin
			nli10iO <= nii00li;
		end
	end
	assign
		wire_nli10il_ENA = (n0O1l & (~ ni1iili));
	event nli10iO_event;
	initial
		#1 ->nli10iO_event;
	always @(nli10iO_event)
		nli10iO <= 1;
	initial
	begin
		nli10lO = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nli10lO <= 0;
		end
		else if  (wire_nli10ll_ENA == 1'b1) 
		begin
			nli10lO <= nl0l1il;
		end
	end
	assign
		wire_nli10ll_ENA = (n0Oll & (~ ni1iili));
	event nli10lO_event;
	initial
		#1 ->nli10lO_event;
	always @(nli10lO_event)
		nli10lO <= 1;
	initial
	begin
		nli10OO = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nli10OO <= 0;
		end
		else if  (wire_nli10Ol_ENA == 1'b1) 
		begin
			nli10OO <= nli10lO;
		end
	end
	assign
		wire_nli10Ol_ENA = (n010O & (~ ni1iili));
	initial
	begin
		nli11lO = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nli11lO <= 0;
		end
		else if  (wire_nli11ll_ENA == 1'b1) 
		begin
			nli11lO <= nii00li;
		end
	end
	assign
		wire_nli11ll_ENA = (n0i0l & (~ ni1iili));
	initial
	begin
		nli11OO = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nli11OO <= 0;
		end
		else if  (wire_nli11Ol_ENA == 1'b1) 
		begin
			nli11OO <= nil10lO;
		end
	end
	assign
		wire_nli11Ol_ENA = (n00Oi & (~ ni1iili));
	initial
	begin
		nli1i0O = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nli1i0O <= 0;
		end
		else if  (wire_nli1i0l_ENA == 1'b1) 
		begin
			nli1i0O <= nli1i1O;
		end
	end
	assign
		wire_nli1i0l_ENA = (n010i & (~ ni1iili));
	event nli1i0O_event;
	initial
		#1 ->nli1i0O_event;
	always @(nli1i0O_event)
		nli1i0O <= 1;
	initial
	begin
		nli1i1O = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nli1i1O <= 0;
		end
		else if  (wire_nli1i1l_ENA == 1'b1) 
		begin
			nli1i1O <= nli10OO;
		end
	end
	assign
		wire_nli1i1l_ENA = (n010l & (~ ni1iili));
	initial
	begin
		nli1iiO = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nli1iiO <= 0;
		end
		else if  (wire_nli1iil_ENA == 1'b1) 
		begin
			nli1iiO <= nli1i0O;
		end
	end
	assign
		wire_nli1iil_ENA = (n011O & (~ ni1iili));
	initial
	begin
		nli1ilO = 0;
	end
	always @ ( posedge clock or  negedge wire_nli1ill_CLRN)
	begin
		if (wire_nli1ill_CLRN == 1'b0) 
		begin
			nli1ilO <= 0;
		end
		else if  (wire_nli1ill_ENA == 1'b1) 
		begin
			nli1ilO <= nli1iiO;
		end
	end
	assign
		wire_nli1ill_ENA = (n1ill & (~ ni1iili)),
		wire_nli1ill_CLRN = ((ni1i10O80 ^ ni1i10O79) & (~ reset));
	initial
	begin
		nli1iOO = 0;
	end
	always @ ( posedge clock or  negedge wire_nli1iOl_CLRN)
	begin
		if (wire_nli1iOl_CLRN == 1'b0) 
		begin
			nli1iOO <= 0;
		end
		else if  (wire_nli1iOl_ENA == 1'b1) 
		begin
			nli1iOO <= ni1i1il;
		end
	end
	assign
		wire_nli1iOl_ENA = (n0O0i & (~ ni1iili)),
		wire_nli1iOl_CLRN = ((ni1i1ii78 ^ ni1i1ii77) & (~ reset));
	event nli1iOO_event;
	initial
		#1 ->nli1iOO_event;
	always @(nli1iOO_event)
		nli1iOO <= 1;
	initial
	begin
		nli1l0i = 0;
		nli1l0l = 0;
		nli1l0O = 0;
		nli1l1l = 0;
		nli1l1O = 0;
		nli1lii = 0;
		nli1lil = 0;
		nli1lli = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nli1l0i <= 0;
			nli1l0l <= 0;
			nli1l0O <= 0;
			nli1l1l <= 0;
			nli1l1O <= 0;
			nli1lii <= 0;
			nli1lil <= 0;
			nli1lli <= 0;
		end
		else if  (ni1i1iO == 1'b1) 
		begin
			nli1l0i <= nl1ii1O;
			nli1l0l <= nl1ii0i;
			nli1l0O <= nl1ii0l;
			nli1l1l <= nl1iili;
			nli1l1O <= nl1ii1l;
			nli1lii <= nl1ii0O;
			nli1lil <= nl1iiii;
			nli1lli <= nl1iiil;
		end
	end
	event nli1l0i_event;
	event nli1l0l_event;
	event nli1l0O_event;
	event nli1l1l_event;
	event nli1l1O_event;
	event nli1lii_event;
	event nli1lil_event;
	event nli1lli_event;
	initial
		#1 ->nli1l0i_event;
	initial
		#1 ->nli1l0l_event;
	initial
		#1 ->nli1l0O_event;
	initial
		#1 ->nli1l1l_event;
	initial
		#1 ->nli1l1O_event;
	initial
		#1 ->nli1lii_event;
	initial
		#1 ->nli1lil_event;
	initial
		#1 ->nli1lli_event;
	always @(nli1l0i_event)
		nli1l0i <= 1;
	always @(nli1l0l_event)
		nli1l0l <= 1;
	always @(nli1l0O_event)
		nli1l0O <= 1;
	always @(nli1l1l_event)
		nli1l1l <= 1;
	always @(nli1l1O_event)
		nli1l1O <= 1;
	always @(nli1lii_event)
		nli1lii <= 1;
	always @(nli1lil_event)
		nli1lil <= 1;
	always @(nli1lli_event)
		nli1lli <= 1;
	initial
	begin
		nli1llO = 0;
		nli1lOi = 0;
		nli1lOl = 0;
		nli1lOO = 0;
		nli1O0l = 0;
		nli1O1i = 0;
		nli1O1l = 0;
		nli1O1O = 0;
	end
	always @ (clock or wire_nli1O0i_PRN or wire_nli1O0i_CLRN)
	begin
		if (wire_nli1O0i_PRN == 1'b0) 
		begin
			nli1llO <= 1;
			nli1lOi <= 1;
			nli1lOl <= 1;
			nli1lOO <= 1;
			nli1O0l <= 1;
			nli1O1i <= 1;
			nli1O1l <= 1;
			nli1O1O <= 1;
		end
		else if  (wire_nli1O0i_CLRN == 1'b0) 
		begin
			nli1llO <= 0;
			nli1lOi <= 0;
			nli1lOl <= 0;
			nli1lOO <= 0;
			nli1O0l <= 0;
			nli1O1i <= 0;
			nli1O1l <= 0;
			nli1O1O <= 0;
		end
		else if  (ni1i1lO == 1'b1) 
		if (clock != nli1O0i_clk_prev && clock == 1'b1) 
		begin
			nli1llO <= nl1il0l;
			nli1lOi <= nl1iilO;
			nli1lOl <= nl1iiOi;
			nli1lOO <= nl1iiOl;
			nli1O0l <= nl1il1O;
			nli1O1i <= nl1iiOO;
			nli1O1l <= nl1il1i;
			nli1O1O <= nl1il1l;
		end
		nli1O0i_clk_prev <= clock;
	end
	assign
		wire_nli1O0i_CLRN = ((ni1i1ll74 ^ ni1i1ll73) & (~ reset)),
		wire_nli1O0i_PRN = (ni1i1li76 ^ ni1i1li75);
	event nli1llO_event;
	event nli1lOi_event;
	event nli1lOl_event;
	event nli1lOO_event;
	event nli1O0l_event;
	event nli1O1i_event;
	event nli1O1l_event;
	event nli1O1O_event;
	initial
		#1 ->nli1llO_event;
	initial
		#1 ->nli1lOi_event;
	initial
		#1 ->nli1lOl_event;
	initial
		#1 ->nli1lOO_event;
	initial
		#1 ->nli1O0l_event;
	initial
		#1 ->nli1O1i_event;
	initial
		#1 ->nli1O1l_event;
	initial
		#1 ->nli1O1O_event;
	always @(nli1llO_event)
		nli1llO <= 1;
	always @(nli1lOi_event)
		nli1lOi <= 1;
	always @(nli1lOl_event)
		nli1lOl <= 1;
	always @(nli1lOO_event)
		nli1lOO <= 1;
	always @(nli1O0l_event)
		nli1O0l <= 1;
	always @(nli1O1i_event)
		nli1O1i <= 1;
	always @(nli1O1l_event)
		nli1O1l <= 1;
	always @(nli1O1O_event)
		nli1O1O <= 1;
	initial
	begin
		nli1Oii = 0;
		nli1Oil = 0;
		nli1OiO = 0;
		nli1Oli = 0;
		nli1Oll = 0;
		nli1OlO = 0;
		nli1OOi = 0;
		nli1OOO = 0;
	end
	always @ (clock or wire_nli1OOl_PRN or wire_nli1OOl_CLRN)
	begin
		if (wire_nli1OOl_PRN == 1'b0) 
		begin
			nli1Oii <= 1;
			nli1Oil <= 1;
			nli1OiO <= 1;
			nli1Oli <= 1;
			nli1Oll <= 1;
			nli1OlO <= 1;
			nli1OOi <= 1;
			nli1OOO <= 1;
		end
		else if  (wire_nli1OOl_CLRN == 1'b0) 
		begin
			nli1Oii <= 0;
			nli1Oil <= 0;
			nli1OiO <= 0;
			nli1Oli <= 0;
			nli1Oll <= 0;
			nli1OlO <= 0;
			nli1OOi <= 0;
			nli1OOO <= 0;
		end
		else if  (ni1i1OO == 1'b1) 
		if (clock != nli1OOl_clk_prev && clock == 1'b1) 
		begin
			nli1Oii <= nl1ilOO;
			nli1Oil <= nl1ilii;
			nli1OiO <= nl1ilil;
			nli1Oli <= nl1iliO;
			nli1Oll <= nl1illi;
			nli1OlO <= nl1illl;
			nli1OOi <= nl1illO;
			nli1OOO <= nl1ilOi;
		end
		nli1OOl_clk_prev <= clock;
	end
	assign
		wire_nli1OOl_CLRN = ((ni1i1Ol70 ^ ni1i1Ol69) & (~ reset)),
		wire_nli1OOl_PRN = (ni1i1Oi72 ^ ni1i1Oi71);
	event nli1Oii_event;
	event nli1Oil_event;
	event nli1OiO_event;
	event nli1Oli_event;
	event nli1Oll_event;
	event nli1OlO_event;
	event nli1OOi_event;
	event nli1OOO_event;
	initial
		#1 ->nli1Oii_event;
	initial
		#1 ->nli1Oil_event;
	initial
		#1 ->nli1OiO_event;
	initial
		#1 ->nli1Oli_event;
	initial
		#1 ->nli1Oll_event;
	initial
		#1 ->nli1OlO_event;
	initial
		#1 ->nli1OOi_event;
	initial
		#1 ->nli1OOO_event;
	always @(nli1Oii_event)
		nli1Oii <= 1;
	always @(nli1Oil_event)
		nli1Oil <= 1;
	always @(nli1OiO_event)
		nli1OiO <= 1;
	always @(nli1Oli_event)
		nli1Oli <= 1;
	always @(nli1Oll_event)
		nli1Oll <= 1;
	always @(nli1OlO_event)
		nli1OlO <= 1;
	always @(nli1OOi_event)
		nli1OOi <= 1;
	always @(nli1OOO_event)
		nli1OOO <= 1;
	initial
	begin
		nlii00l = 0;
		nlii01i = 0;
		nlii01l = 0;
		nlii01O = 0;
	end
	always @ ( posedge clock or  negedge wire_nlii00i_CLRN)
	begin
		if (wire_nlii00i_CLRN == 1'b0) 
		begin
			nlii00l <= 0;
			nlii01i <= 0;
			nlii01l <= 0;
			nlii01O <= 0;
		end
		else if  (ni1ii0i == 1'b1) 
		begin
			nlii00l <= nii10il;
			nlii01i <= nii100l;
			nlii01l <= nii100O;
			nlii01O <= nii10ii;
		end
	end
	assign
		wire_nlii00i_CLRN = ((ni1ii1O48 ^ ni1ii1O47) & (~ reset));
	event nlii00l_event;
	event nlii01i_event;
	event nlii01l_event;
	event nlii01O_event;
	initial
		#1 ->nlii00l_event;
	initial
		#1 ->nlii01i_event;
	initial
		#1 ->nlii01l_event;
	initial
		#1 ->nlii01O_event;
	always @(nlii00l_event)
		nlii00l <= 1;
	always @(nlii01i_event)
		nlii01i <= 1;
	always @(nlii01l_event)
		nlii01l <= 1;
	always @(nlii01O_event)
		nlii01O <= 1;
	initial
	begin
		nlii0ii = 0;
		nlii0il = 0;
		nlii0iO = 0;
		nlii0ll = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nlii0ii <= 0;
			nlii0il <= 0;
			nlii0iO <= 0;
			nlii0ll <= 0;
		end
		else if  (ni1ii0l == 1'b1) 
		begin
			nlii0ii <= nii10Oi;
			nlii0il <= nii10Ol;
			nlii0iO <= nii10OO;
			nlii0ll <= nii1i1i;
		end
	end
	event nlii0ii_event;
	event nlii0il_event;
	event nlii0iO_event;
	event nlii0ll_event;
	initial
		#1 ->nlii0ii_event;
	initial
		#1 ->nlii0il_event;
	initial
		#1 ->nlii0iO_event;
	initial
		#1 ->nlii0ll_event;
	always @(nlii0ii_event)
		nlii0ii <= 1;
	always @(nlii0il_event)
		nlii0il <= 1;
	always @(nlii0iO_event)
		nlii0iO <= 1;
	always @(nlii0ll_event)
		nlii0ll <= 1;
	initial
	begin
		nli0O0i = 0;
		nli0O0l = 0;
		nli0O0O = 0;
		nli0O1l = 0;
		nli0O1O = 0;
		nli0Oii = 0;
		nli0Oil = 0;
		nli0OiO = 0;
		nli0Oli = 0;
		nli0Oll = 0;
		nli0OlO = 0;
		nli0OOi = 0;
		nli0OOl = 0;
		nli0OOO = 0;
		nlii10i = 0;
		nlii10l = 0;
		nlii10O = 0;
		nlii11i = 0;
		nlii11l = 0;
		nlii11O = 0;
		nlii1ii = 0;
		nlii1il = 0;
		nlii1iO = 0;
		nlii1ll = 0;
	end
	always @ (clock or wire_nlii1li_PRN or reset)
	begin
		if (wire_nlii1li_PRN == 1'b0) 
		begin
			nli0O0i <= 1;
			nli0O0l <= 1;
			nli0O0O <= 1;
			nli0O1l <= 1;
			nli0O1O <= 1;
			nli0Oii <= 1;
			nli0Oil <= 1;
			nli0OiO <= 1;
			nli0Oli <= 1;
			nli0Oll <= 1;
			nli0OlO <= 1;
			nli0OOi <= 1;
			nli0OOl <= 1;
			nli0OOO <= 1;
			nlii10i <= 1;
			nlii10l <= 1;
			nlii10O <= 1;
			nlii11i <= 1;
			nlii11l <= 1;
			nlii11O <= 1;
			nlii1ii <= 1;
			nlii1il <= 1;
			nlii1iO <= 1;
			nlii1ll <= 1;
		end
		else if  (reset == 1'b1) 
		begin
			nli0O0i <= 0;
			nli0O0l <= 0;
			nli0O0O <= 0;
			nli0O1l <= 0;
			nli0O1O <= 0;
			nli0Oii <= 0;
			nli0Oil <= 0;
			nli0OiO <= 0;
			nli0Oli <= 0;
			nli0Oll <= 0;
			nli0OlO <= 0;
			nli0OOi <= 0;
			nli0OOl <= 0;
			nli0OOO <= 0;
			nlii10i <= 0;
			nlii10l <= 0;
			nlii10O <= 0;
			nlii11i <= 0;
			nlii11l <= 0;
			nlii11O <= 0;
			nlii1ii <= 0;
			nlii1il <= 0;
			nlii1iO <= 0;
			nlii1ll <= 0;
		end
		else if  (ni1ii1l == 1'b1) 
		if (clock != nlii1li_clk_prev && clock == 1'b1) 
		begin
			nli0O0i <= nii11Ol;
			nli0O0l <= nii11OO;
			nli0O0O <= nii101i;
			nli0O1l <= nii11lO;
			nli0O1O <= nii11Oi;
			nli0Oii <= nii101l;
			nli0Oil <= nii101O;
			nli0OiO <= nii100i;
			nli0Oli <= nii100l;
			nli0Oll <= nii100O;
			nli0OlO <= nii10ii;
			nli0OOi <= nii10il;
			nli0OOl <= nii10iO;
			nli0OOO <= nii10li;
			nlii10i <= nii10Ol;
			nlii10l <= nii10OO;
			nlii10O <= nii1i1i;
			nlii11i <= nii10ll;
			nlii11l <= nii10lO;
			nlii11O <= nii10Oi;
			nlii1ii <= nii1i1l;
			nlii1il <= nii1i1O;
			nlii1iO <= nii1i0i;
			nlii1ll <= nii1i0l;
		end
		nlii1li_clk_prev <= clock;
	end
	assign
		wire_nlii1li_PRN = (ni1ii1i50 ^ ni1ii1i49);
	event nli0O0i_event;
	event nli0O0l_event;
	event nli0O0O_event;
	event nli0O1l_event;
	event nli0O1O_event;
	event nli0Oii_event;
	event nli0Oil_event;
	event nli0OiO_event;
	event nli0Oli_event;
	event nli0Oll_event;
	event nli0OlO_event;
	event nli0OOi_event;
	event nli0OOl_event;
	event nli0OOO_event;
	event nlii10i_event;
	event nlii10l_event;
	event nlii10O_event;
	event nlii11i_event;
	event nlii11l_event;
	event nlii11O_event;
	event nlii1ii_event;
	event nlii1il_event;
	event nlii1iO_event;
	event nlii1ll_event;
	initial
		#1 ->nli0O0i_event;
	initial
		#1 ->nli0O0l_event;
	initial
		#1 ->nli0O0O_event;
	initial
		#1 ->nli0O1l_event;
	initial
		#1 ->nli0O1O_event;
	initial
		#1 ->nli0Oii_event;
	initial
		#1 ->nli0Oil_event;
	initial
		#1 ->nli0OiO_event;
	initial
		#1 ->nli0Oli_event;
	initial
		#1 ->nli0Oll_event;
	initial
		#1 ->nli0OlO_event;
	initial
		#1 ->nli0OOi_event;
	initial
		#1 ->nli0OOl_event;
	initial
		#1 ->nli0OOO_event;
	initial
		#1 ->nlii10i_event;
	initial
		#1 ->nlii10l_event;
	initial
		#1 ->nlii10O_event;
	initial
		#1 ->nlii11i_event;
	initial
		#1 ->nlii11l_event;
	initial
		#1 ->nlii11O_event;
	initial
		#1 ->nlii1ii_event;
	initial
		#1 ->nlii1il_event;
	initial
		#1 ->nlii1iO_event;
	initial
		#1 ->nlii1ll_event;
	always @(nli0O0i_event)
		nli0O0i <= 1;
	always @(nli0O0l_event)
		nli0O0l <= 1;
	always @(nli0O0O_event)
		nli0O0O <= 1;
	always @(nli0O1l_event)
		nli0O1l <= 1;
	always @(nli0O1O_event)
		nli0O1O <= 1;
	always @(nli0Oii_event)
		nli0Oii <= 1;
	always @(nli0Oil_event)
		nli0Oil <= 1;
	always @(nli0OiO_event)
		nli0OiO <= 1;
	always @(nli0Oli_event)
		nli0Oli <= 1;
	always @(nli0Oll_event)
		nli0Oll <= 1;
	always @(nli0OlO_event)
		nli0OlO <= 1;
	always @(nli0OOi_event)
		nli0OOi <= 1;
	always @(nli0OOl_event)
		nli0OOl <= 1;
	always @(nli0OOO_event)
		nli0OOO <= 1;
	always @(nlii10i_event)
		nlii10i <= 1;
	always @(nlii10l_event)
		nlii10l <= 1;
	always @(nlii10O_event)
		nlii10O <= 1;
	always @(nlii11i_event)
		nlii11i <= 1;
	always @(nlii11l_event)
		nlii11l <= 1;
	always @(nlii11O_event)
		nlii11O <= 1;
	always @(nlii1ii_event)
		nlii1ii <= 1;
	always @(nlii1il_event)
		nlii1il <= 1;
	always @(nlii1iO_event)
		nlii1iO <= 1;
	always @(nlii1ll_event)
		nlii1ll <= 1;
	initial
	begin
		nlii1Ol = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nlii1Ol <= 0;
		end
		else if  (wire_nlii1Oi_ENA == 1'b1) 
		begin
			nlii1Ol <= nl0l0Oi;
		end
	end
	assign
		wire_nlii1Oi_ENA = (n111l & (~ ni1iiii));
	initial
	begin
		nlii0Oi = 0;
		nlii0Ol = 0;
		nlii0OO = 0;
		nliii1l = 0;
	end
	always @ ( posedge clock or  posedge reset)
	begin
		if (reset == 1'b1) 
		begin
			nlii0Oi <= 0;
			nlii0Ol <= 0;
			nlii0OO <= 0;
			nliii1l <= 0;
		end
		else if  (ni1ii0O == 1'b1) 
		begin
			nlii0Oi <= nlii0ii;
			nlii0Ol <= nlii0il;
			nlii0OO <= nlii0iO;
			nliii1l <= nlii0ll;
		end
	end
	initial
	begin
		ni0000i = 0;
		ni0000O = 0;
		ni0001l = 0;
		ni000ii = 0;
		ni000iO = 0;
		ni000ll = 0;
		ni000Oi = 0;
		ni000Ol = 0;
		ni000OO = 0;
		ni0010i = 0;
		ni0010l = 0;
		ni0010O = 0;
		ni0011i = 0;
		ni0011O = 0;
		ni001il = 0;
		ni001iO = 0;
		ni001li = 0;
		ni001lO = 0;
		ni001Oi = 0;
		ni001OO = 0;
		ni00i0i = 0;
		ni00i0l = 0;
		ni00i1i = 0;
		ni00i1O = 0;
		ni00iii = 0;
		ni00iil = 0;
		ni00ili = 0;
		ni00ilO = 0;
		ni00iOl = 0;
		ni00l0i = 0;
		ni00l0O = 0;
		ni00l1i = 0;
		ni00l1l = 0;
		ni00lil = 0;
		ni00liO = 0;
		ni00lli = 0;
		ni00lll = 0;
		ni00lOi = 0;
		ni00lOl = 0;
		ni00lOO = 0;
		ni00O0l = 0;
		ni00O1l = 0;
		ni00O1O = 0;
		ni00Oii = 0;
		ni0100O = 0;
		ni01Oll = 0;
		ni01OlO = 0;
		ni01OOl = 0;
		ni0il1O = 0;
		nl001li = 0;
		nl001ll = 0;
		nl01O0l = 0;
		nl01O0O = 0;
		nllOOO = 0;
		nlO1Oi = 0;
	end
	always @ (clock or reset or wire_nlO1lO_CLRN)
	begin
		if (reset == 1'b1) 
		begin
			ni0000i <= 1;
			ni0000O <= 1;
			ni0001l <= 1;
			ni000ii <= 1;
			ni000iO <= 1;
			ni000ll <= 1;
			ni000Oi <= 1;
			ni000Ol <= 1;
			ni000OO <= 1;
			ni0010i <= 1;
			ni0010l <= 1;
			ni0010O <= 1;
			ni0011i <= 1;
			ni0011O <= 1;
			ni001il <= 1;
			ni001iO <= 1;
			ni001li <= 1;
			ni001lO <= 1;
			ni001Oi <= 1;
			ni001OO <= 1;
			ni00i0i <= 1;
			ni00i0l <= 1;
			ni00i1i <= 1;
			ni00i1O <= 1;
			ni00iii <= 1;
			ni00iil <= 1;
			ni00ili <= 1;
			ni00ilO <= 1;
			ni00iOl <= 1;
			ni00l0i <= 1;
			ni00l0O <= 1;
			ni00l1i <= 1;
			ni00l1l <= 1;
			ni00lil <= 1;
			ni00liO <= 1;
			ni00lli <= 1;
			ni00lll <= 1;
			ni00lOi <= 1;
			ni00lOl <= 1;
			ni00lOO <= 1;
			ni00O0l <= 1;
			ni00O1l <= 1;
			ni00O1O <= 1;
			ni00Oii <= 1;
			ni0100O <= 1;
			ni01Oll <= 1;
			ni01OlO <= 1;
			ni01OOl <= 1;
			ni0il1O <= 1;
			nl001li <= 1;
			nl001ll <= 1;
			nl01O0l <= 1;
			nl01O0O <= 1;
			nllOOO <= 1;
			nlO1Oi <= 1;
		end
		else if  (wire_nlO1lO_CLRN == 1'b0) 
		begin
			ni0000i <= 0;
			ni0000O <= 0;
			ni0001l <= 0;
			ni000ii <= 0;
			ni000iO <= 0;
			ni000ll <= 0;
			ni000Oi <= 0;
			ni000Ol <= 0;
			ni000OO <= 0;
			ni0010i <= 0;
			ni0010l <= 0;
			ni0010O <= 0;
			ni0011i <= 0;
			ni0011O <= 0;
			ni001il <= 0;
			ni001iO <= 0;
			ni001li <= 0;
			ni001lO <= 0;
			ni001Oi <= 0;
			ni001OO <= 0;
			ni00i0i <= 0;
			ni00i0l <= 0;
			ni00i1i <= 0;
			ni00i1O <= 0;
			ni00iii <= 0;
			ni00iil <= 0;
			ni00ili <= 0;
			ni00ilO <= 0;
			ni00iOl <= 0;
			ni00l0i <= 0;
			ni00l0O <= 0;
			ni00l1i <= 0;
			ni00l1l <= 0;
			ni00lil <= 0;
			ni00liO <= 0;
			ni00lli <= 0;
			ni00lll <= 0;
			ni00lOi <= 0;
			ni00lOl <= 0;
			ni00lOO <= 0;
			ni00O0l <= 0;
			ni00O1l <= 0;
			ni00O1O <= 0;
			ni00Oii <= 0;
			ni0100O <= 0;
			ni01Oll <= 0;
			ni01OlO <= 0;
			ni01OOl <= 0;
			ni0il1O <= 0;
			nl001li <= 0;
			nl001ll <= 0;
			nl01O0l <= 0;
			nl01O0O <= 0;
			nllOOO <= 0;
			nlO1Oi <= 0;
		end
		else 
		if (clock != nlO1lO_clk_prev && clock == 1'b1) 
		begin
			ni0000i <= wire_ni0il0i_dataout;
			ni0000O <= wire_ni0il0O_dataout;
			ni0001l <= wire_ni0ll0O_dataout;
			ni000ii <= wire_ni0ilii_dataout;
			ni000iO <= wire_ni0iliO_dataout;
			ni000ll <= wire_ni0illl_dataout;
			ni000Oi <= wire_ni0ilOi_dataout;
			ni000Ol <= wire_ni0ilOl_dataout;
			ni000OO <= wire_ni0ilOO_dataout;
			ni0010i <= wire_ni0liil_dataout;
			ni0010l <= wire_ni0liiO_dataout;
			ni0010O <= wire_ni0lili_dataout;
			ni0011i <= wire_ni0li0l_dataout;
			ni0011O <= wire_ni0liii_dataout;
			ni001il <= wire_ni0lilO_dataout;
			ni001iO <= wire_ni0liOi_dataout;
			ni001li <= wire_ni0liOl_dataout;
			ni001lO <= wire_ni0ll1i_dataout;
			ni001Oi <= wire_ni0ll1l_dataout;
			ni001OO <= wire_ni0ll0i_dataout;
			ni00i0i <= wire_ni0iO0i_dataout;
			ni00i0l <= wire_ni0iO0l_dataout;
			ni00i1i <= wire_ni0iO1i_dataout;
			ni00i1O <= wire_ni0iO1O_dataout;
			ni00iii <= wire_ni0iOii_dataout;
			ni00iil <= wire_ni0iOil_dataout;
			ni00ili <= wire_ni0iOli_dataout;
			ni00ilO <= wire_ni0iOlO_dataout;
			ni00iOl <= wire_ni00OiO_dataout;
			ni00l0i <= wire_ni00OOl_dataout;
			ni00l0O <= wire_ni0i11i_dataout;
			ni00l1i <= wire_ni00Oll_dataout;
			ni00l1l <= wire_ni00OlO_dataout;
			ni00lil <= wire_ni0i11O_dataout;
			ni00liO <= wire_ni0i10i_dataout;
			ni00lli <= wire_ni0i10l_dataout;
			ni00lll <= wire_ni0i10O_dataout;
			ni00lOi <= wire_ni0i1il_dataout;
			ni00lOl <= wire_ni0i1iO_dataout;
			ni00lOO <= wire_ni0i1li_dataout;
			ni00O0l <= wire_ni0i1OO_dataout;
			ni00O1l <= wire_ni0i1lO_dataout;
			ni00O1O <= wire_ni0i1Oi_dataout;
			ni00Oii <= wire_ni0i01l_dataout;
			ni0100O <= wire_ni010lO_dataout;
			ni01Oll <= wire_ni0l0OO_dataout;
			ni01OlO <= wire_ni0li1i_dataout;
			ni01OOl <= wire_ni0li1O_dataout;
			ni0il1O <= wire_ni0l0Oi_dataout;
			nl001li <= nl001ll;
			nl001ll <= ni10O1l;
			nl01O0l <= nl01O0O;
			nl01O0O <= ni10O1l;
			nllOOO <= nl01O0O;
			nlO1Oi <= nl001ll;
		end
		nlO1lO_clk_prev <= clock;
	end
	assign
		wire_nlO1lO_CLRN = (ni1iill46 ^ ni1iill45);
	event ni0000i_event;
	event ni0000O_event;
	event ni0001l_event;
	event ni000ii_event;
	event ni000iO_event;
	event ni000ll_event;
	event ni000Oi_event;
	event ni000Ol_event;
	event ni000OO_event;
	event ni0010i_event;
	event ni0010l_event;
	event ni0010O_event;
	event ni0011i_event;
	event ni0011O_event;
	event ni001il_event;
	event ni001iO_event;
	event ni001li_event;
	event ni001lO_event;
	event ni001Oi_event;
	event ni001OO_event;
	event ni00i0i_event;
	event ni00i0l_event;
	event ni00i1i_event;
	event ni00i1O_event;
	event ni00iii_event;
	event ni00iil_event;
	event ni00ili_event;
	event ni00ilO_event;
	event ni00iOl_event;
	event ni00l0i_event;
	event ni00l0O_event;
	event ni00l1i_event;
	event ni00l1l_event;
	event ni00lil_event;
	event ni00liO_event;
	event ni00lli_event;
	event ni00lll_event;
	event ni00lOi_event;
	event ni00lOl_event;
	event ni00lOO_event;
	event ni00O0l_event;
	event ni00O1l_event;
	event ni00O1O_event;
	event ni00Oii_event;
	event ni0100O_event;
	event ni01Oll_event;
	event ni01OlO_event;
	event ni01OOl_event;
	event ni0il1O_event;
	event nl001li_event;
	event nl001ll_event;
	event nl01O0l_event;
	event nl01O0O_event;
	event nllOOO_event;
	event nlO1Oi_event;
	initial
		#1 ->ni0000i_event;
	initial
		#1 ->ni0000O_event;
	initial
		#1 ->ni0001l_event;
	initial
		#1 ->ni000ii_event;
	initial
		#1 ->ni000iO_event;
	initial
		#1 ->ni000ll_event;
	initial
		#1 ->ni000Oi_event;
	initial
		#1 ->ni000Ol_event;
	initial
		#1 ->ni000OO_event;
	initial
		#1 ->ni0010i_event;
	initial
		#1 ->ni0010l_event;
	initial
		#1 ->ni0010O_event;
	initial
		#1 ->ni0011i_event;
	initial
		#1 ->ni0011O_event;
	initial
		#1 ->ni001il_event;
	initial
		#1 ->ni001iO_event;
	initial
		#1 ->ni001li_event;
	initial
		#1 ->ni001lO_event;
	initial
		#1 ->ni001Oi_event;
	initial
		#1 ->ni001OO_event;
	initial
		#1 ->ni00i0i_event;
	initial
		#1 ->ni00i0l_event;
	initial
		#1 ->ni00i1i_event;
	initial
		#1 ->ni00i1O_event;
	initial
		#1 ->ni00iii_event;
	initial
		#1 ->ni00iil_event;
	initial
		#1 ->ni00ili_event;
	initial
		#1 ->ni00ilO_event;
	initial
		#1 ->ni00iOl_event;
	initial
		#1 ->ni00l0i_event;
	initial
		#1 ->ni00l0O_event;
	initial
		#1 ->ni00l1i_event;
	initial
		#1 ->ni00l1l_event;
	initial
		#1 ->ni00lil_event;
	initial
		#1 ->ni00liO_event;
	initial
		#1 ->ni00lli_event;
	initial
		#1 ->ni00lll_event;
	initial
		#1 ->ni00lOi_event;
	initial
		#1 ->ni00lOl_event;
	initial
		#1 ->ni00lOO_event;
	initial
		#1 ->ni00O0l_event;
	initial
		#1 ->ni00O1l_event;
	initial
		#1 ->ni00O1O_event;
	initial
		#1 ->ni00Oii_event;
	initial
		#1 ->ni0100O_event;
	initial
		#1 ->ni01Oll_event;
	initial
		#1 ->ni01OlO_event;
	initial
		#1 ->ni01OOl_event;
	initial
		#1 ->ni0il1O_event;
	initial
		#1 ->nl001li_event;
	initial
		#1 ->nl001ll_event;
	initial
		#1 ->nl01O0l_event;
	initial
		#1 ->nl01O0O_event;
	initial
		#1 ->nllOOO_event;
	initial
		#1 ->nlO1Oi_event;
	always @(ni0000i_event)
		ni0000i <= 1;
	always @(ni0000O_event)
		ni0000O <= 1;
	always @(ni0001l_event)
		ni0001l <= 1;
	always @(ni000ii_event)
		ni000ii <= 1;
	always @(ni000iO_event)
		ni000iO <= 1;
	always @(ni000ll_event)
		ni000ll <= 1;
	always @(ni000Oi_event)
		ni000Oi <= 1;
	always @(ni000Ol_event)
		ni000Ol <= 1;
	always @(ni000OO_event)
		ni000OO <= 1;
	always @(ni0010i_event)
		ni0010i <= 1;
	always @(ni0010l_event)
		ni0010l <= 1;
	always @(ni0010O_event)
		ni0010O <= 1;
	always @(ni0011i_event)
		ni0011i <= 1;
	always @(ni0011O_event)
		ni0011O <= 1;
	always @(ni001il_event)
		ni001il <= 1;
	always @(ni001iO_event)
		ni001iO <= 1;
	always @(ni001li_event)
		ni001li <= 1;
	always @(ni001lO_event)
		ni001lO <= 1;
	always @(ni001Oi_event)
		ni001Oi <= 1;
	always @(ni001OO_event)
		ni001OO <= 1;
	always @(ni00i0i_event)
		ni00i0i <= 1;
	always @(ni00i0l_event)
		ni00i0l <= 1;
	always @(ni00i1i_event)
		ni00i1i <= 1;
	always @(ni00i1O_event)
		ni00i1O <= 1;
	always @(ni00iii_event)
		ni00iii <= 1;
	always @(ni00iil_event)
		ni00iil <= 1;
	always @(ni00ili_event)
		ni00ili <= 1;
	always @(ni00ilO_event)
		ni00ilO <= 1;
	always @(ni00iOl_event)
		ni00iOl <= 1;
	always @(ni00l0i_event)
		ni00l0i <= 1;
	always @(ni00l0O_event)
		ni00l0O <= 1;
	always @(ni00l1i_event)
		ni00l1i <= 1;
	always @(ni00l1l_event)
		ni00l1l <= 1;
	always @(ni00lil_event)
		ni00lil <= 1;
	always @(ni00liO_event)
		ni00liO <= 1;
	always @(ni00lli_event)
		ni00lli <= 1;
	always @(ni00lll_event)
		ni00lll <= 1;
	always @(ni00lOi_event)
		ni00lOi <= 1;
	always @(ni00lOl_event)
		ni00lOl <= 1;
	always @(ni00lOO_event)
		ni00lOO <= 1;
	always @(ni00O0l_event)
		ni00O0l <= 1;
	always @(ni00O1l_event)
		ni00O1l <= 1;
	always @(ni00O1O_event)
		ni00O1O <= 1;
	always @(ni00Oii_event)
		ni00Oii <= 1;
	always @(ni0100O_event)
		ni0100O <= 1;
	always @(ni01Oll_event)
		ni01Oll <= 1;
	always @(ni01OlO_event)
		ni01OlO <= 1;
	always @(ni01OOl_event)
		ni01OOl <= 1;
	always @(ni0il1O_event)
		ni0il1O <= 1;
	always @(nl001li_event)
		nl001li <= 1;
	always @(nl001ll_event)
		nl001ll <= 1;
	always @(nl01O0l_event)
		nl01O0l <= 1;
	always @(nl01O0O_event)
		nl01O0O <= 1;
	always @(nllOOO_event)
		nllOOO <= 1;
	always @(nlO1Oi_event)
		nlO1Oi <= 1;
	lpm_counter   nl001iO
	( 
	.aset(reset),
	.clk_en(ni1iiOO),
	.clock(clock),
	.cout(),
	.data({wire_nlO1ll_o, wire_nlO1li_o, wire_nlO1iO_o, wire_nlO1il_o, n110i, wire_nlO1ii_o, wire_nlO10O_o}),
	.q(wire_nl001iO_q),
	.sload(((~ ni1iiii) & wire_nl0010O_o)),
	.aclr(),
	.aload(),
	.cin(),
	.cnt_en(),
	.sclr(),
	.sset(),
	.updown()
	);
	defparam
		nl001iO.lpm_avalue = "0",
		nl001iO.lpm_direction = "UP",
		nl001iO.lpm_modulus = 0,
		nl001iO.lpm_port_updown = "PORT_CONNECTIVITY",
		nl001iO.lpm_width = 7;
	lpm_counter   nl01O0i
	( 
	.aset(reset),
	.clk_en(ni1il1l),
	.clock(clock),
	.cout(),
	.data({n0Oll, n001O, n00ii, n001l, n0Oil, n001i, n01OO, n01Ol}),
	.q(wire_nl01O0i_q),
	.sload(((~ ni1iili) & wire_nl01lii_o)),
	.aclr(),
	.aload(),
	.cin(),
	.cnt_en(),
	.sclr(),
	.sset(),
	.updown()
	);
	defparam
		nl01O0i.lpm_avalue = "0",
		nl01O0i.lpm_direction = "UP",
		nl01O0i.lpm_modulus = 0,
		nl01O0i.lpm_port_updown = "PORT_CONNECTIVITY",
		nl01O0i.lpm_width = 8;
	assign		wire_ni00OiO_dataout = (n0OOlOO === 1'b1) ? wire_ni1l11O_dataout : wire_ni0i00i_dataout;
	assign		wire_ni00Oli_dataout = (n0OOlOO === 1'b1) ? wire_ni1l10i_dataout : wire_ni0i00l_dataout;
	assign		wire_ni00Oll_dataout = (n0OOlOO === 1'b1) ? wire_ni1l10l_dataout : wire_ni0i00O_dataout;
	assign		wire_ni00OlO_dataout = (n0OOlOO === 1'b1) ? wire_ni1l10O_dataout : wire_ni0i0ii_dataout;
	assign		wire_ni00OOi_dataout = (n0OOlOO === 1'b1) ? wire_ni1l1ii_dataout : wire_ni0i0il_dataout;
	assign		wire_ni00OOl_dataout = (n0OOlOO === 1'b1) ? wire_ni1l1il_dataout : wire_ni0i0iO_dataout;
	assign		wire_ni00OOO_dataout = (n0OOlOO === 1'b1) ? wire_ni1l1iO_dataout : wire_ni0i0li_dataout;
	assign		wire_ni010il_dataout = (n0OOlli === 1'b1) ? wire_ni01i1l_o[1] : wire_ni010li_dataout;
	assign		wire_ni010iO_dataout = (n0OOlli === 1'b1) ? wire_ni01i1l_o[2] : wire_ni010ll_dataout;
	assign		wire_ni010li_dataout = (n0OOliO === 1'b1) ? wire_ni010Ol_o[0] : ni01i1O;
	assign		wire_ni010ll_dataout = (n0OOliO === 1'b1) ? wire_ni010Ol_o[1] : ni0100l;
	assign		wire_ni010lO_dataout = (n0OOlli === 1'b1) ? wire_ni01i0i_dataout : wire_ni010Oi_dataout;
	and(wire_ni010Oi_dataout, ni0100O, ~(n0OOliO));
	and(wire_ni0111i_dataout, nl10l1O, n0OOiOO);
	and(wire_ni0111l_dataout, nli11OO, n0OOiOO);
	or(wire_ni01i0i_dataout, ni0100O, (ni01i1O & (~ ni0100l)));
	assign		wire_ni01iiO_dataout = (n0OOllO === 1'b1) ? wire_ni01l0i_o[1] : wire_ni01ill_dataout;
	assign		wire_ni01ili_dataout = (n0OOllO === 1'b1) ? wire_ni01l0i_o[2] : wire_ni01ilO_dataout;
	assign		wire_ni01ill_dataout = (n0OOlll === 1'b1) ? wire_ni01iOO_o[0] : ni010ii;
	assign		wire_ni01ilO_dataout = (n0OOlll === 1'b1) ? wire_ni01iOO_o[1] : ni01iii;
	and(wire_ni01iOi_dataout, wire_ni01iOl_dataout, ~(n0OOllO));
	assign		wire_ni01iOl_dataout = (n0OOlll === 1'b1) ? wire_ni01l1i_dataout : ni01iil;
	or(wire_ni01l1i_dataout, ni01iil, (ni01iii & (~ ni010ii)));
	assign		wire_ni01lll_dataout = (n0OOlOl === 1'b1) ? wire_ni01O1O_o[1] : wire_ni01lOi_dataout;
	assign		wire_ni01llO_dataout = (n0OOlOl === 1'b1) ? wire_ni01O1O_o[2] : wire_ni01lOl_dataout;
	assign		wire_ni01lOi_dataout = (n0OOlOi === 1'b1) ? wire_ni01lOO_o[0] : ni01liO;
	assign		wire_ni01lOl_dataout = (n0OOlOi === 1'b1) ? wire_ni01lOO_o[1] : ni01lli;
	or(wire_ni0i00i_dataout, ni00iOl, n0OOO0l);
	and(wire_ni0i00l_dataout, ni00iOO, ~(n0OOO0l));
	or(wire_ni0i00O_dataout, ni00l1i, n0OOO0l);
	assign		wire_ni0i01i_dataout = (n0OOlOO === 1'b1) ? wire_ni1l0li_dataout : wire_ni0iill_dataout;
	assign		wire_ni0i01l_dataout = (n0OOlOO === 1'b1) ? wire_ni1l0ll_dataout : wire_ni0iilO_dataout;
	assign		wire_ni0i01O_dataout = (n0OOlOO === 1'b1) ? wire_ni1l0lO_dataout : wire_ni0iiOi_dataout;
	or(wire_ni0i0ii_dataout, ni00l1l, n0OOO0l);
	and(wire_ni0i0il_dataout, ni00l1O, ~(n0OOO0l));
	or(wire_ni0i0iO_dataout, ni00l0i, n0OOO0l);
	and(wire_ni0i0li_dataout, ni00l0l, ~(n0OOO0l));
	or(wire_ni0i0ll_dataout, ni00l0O, n0OOO0l);
	and(wire_ni0i0lO_dataout, ni00lii, ~(n0OOO0l));
	or(wire_ni0i0Oi_dataout, ni00lil, n0OOO0l);
	or(wire_ni0i0Ol_dataout, ni00liO, n0OOO0l);
	or(wire_ni0i0OO_dataout, ni00lli, n0OOO0l);
	assign		wire_ni0i10i_dataout = (n0OOlOO === 1'b1) ? wire_ni1l1Oi_dataout : wire_ni0i0Ol_dataout;
	assign		wire_ni0i10l_dataout = (n0OOlOO === 1'b1) ? wire_ni1l1Ol_dataout : wire_ni0i0OO_dataout;
	assign		wire_ni0i10O_dataout = (n0OOlOO === 1'b1) ? wire_ni1l1OO_dataout : wire_ni0ii1i_dataout;
	assign		wire_ni0i11i_dataout = (n0OOlOO === 1'b1) ? wire_ni1l1li_dataout : wire_ni0i0ll_dataout;
	assign		wire_ni0i11l_dataout = (n0OOlOO === 1'b1) ? wire_ni1l1ll_dataout : wire_ni0i0lO_dataout;
	assign		wire_ni0i11O_dataout = (n0OOlOO === 1'b1) ? wire_ni1l1lO_dataout : wire_ni0i0Oi_dataout;
	assign		wire_ni0i1ii_dataout = (n0OOlOO === 1'b1) ? wire_ni1l01i_dataout : wire_ni0ii1l_dataout;
	assign		wire_ni0i1il_dataout = (n0OOlOO === 1'b1) ? wire_ni1l01l_dataout : wire_ni0ii1O_dataout;
	assign		wire_ni0i1iO_dataout = (n0OOlOO === 1'b1) ? wire_ni1l01O_dataout : wire_ni0ii0i_dataout;
	assign		wire_ni0i1li_dataout = (n0OOlOO === 1'b1) ? wire_ni1l00i_dataout : wire_ni0ii0l_dataout;
	assign		wire_ni0i1ll_dataout = (n0OOlOO === 1'b1) ? wire_ni1l00l_dataout : wire_ni0ii0O_dataout;
	assign		wire_ni0i1lO_dataout = (n0OOlOO === 1'b1) ? wire_ni1l00O_dataout : wire_ni0iiii_dataout;
	assign		wire_ni0i1Oi_dataout = (n0OOlOO === 1'b1) ? wire_ni1l0ii_dataout : wire_ni0iiil_dataout;
	assign		wire_ni0i1Ol_dataout = (n0OOlOO === 1'b1) ? wire_ni1l0il_dataout : wire_ni0iiiO_dataout;
	assign		wire_ni0i1OO_dataout = (n0OOlOO === 1'b1) ? wire_ni1l0iO_dataout : wire_ni0iili_dataout;
	or(wire_ni0ii0i_dataout, ni00lOl, n0OOO0l);
	or(wire_ni0ii0l_dataout, ni00lOO, n0OOO0l);
	and(wire_ni0ii0O_dataout, ni00O1i, ~(n0OOO0l));
	or(wire_ni0ii1i_dataout, ni00lll, n0OOO0l);
	and(wire_ni0ii1l_dataout, ni00llO, ~(n0OOO0l));
	or(wire_ni0ii1O_dataout, ni00lOi, n0OOO0l);
	or(wire_ni0iiii_dataout, ni00O1l, n0OOO0l);
	or(wire_ni0iiil_dataout, ni00O1O, n0OOO0l);
	and(wire_ni0iiiO_dataout, ni00O0i, ~(n0OOO0l));
	or(wire_ni0iili_dataout, ni00O0l, n0OOO0l);
	and(wire_ni0iill_dataout, ni00O0O, ~(n0OOO0l));
	or(wire_ni0iilO_dataout, ni00Oii, n0OOO0l);
	and(wire_ni0iiOi_dataout, ni00Oil, ~(n0OOO0l));
	assign		wire_ni0il0i_dataout = (n0OOO1i === 1'b1) ? wire_ni1l11O_dataout : wire_ni0iOOl_dataout;
	assign		wire_ni0il0l_dataout = (n0OOO1i === 1'b1) ? wire_ni1l10i_dataout : wire_ni0iOOO_dataout;
	assign		wire_ni0il0O_dataout = (n0OOO1i === 1'b1) ? wire_ni1l10l_dataout : wire_ni0l11i_dataout;
	assign		wire_ni0ilii_dataout = (n0OOO1i === 1'b1) ? wire_ni1l10O_dataout : wire_ni0l11l_dataout;
	assign		wire_ni0ilil_dataout = (n0OOO1i === 1'b1) ? wire_ni1l1ii_dataout : wire_ni0l11O_dataout;
	assign		wire_ni0iliO_dataout = (n0OOO1i === 1'b1) ? wire_ni1l1il_dataout : wire_ni0l10i_dataout;
	assign		wire_ni0illi_dataout = (n0OOO1i === 1'b1) ? wire_ni1l1iO_dataout : wire_ni0l10l_dataout;
	assign		wire_ni0illl_dataout = (n0OOO1i === 1'b1) ? wire_ni1l1li_dataout : wire_ni0l10O_dataout;
	assign		wire_ni0illO_dataout = (n0OOO1i === 1'b1) ? wire_ni1l1ll_dataout : wire_ni0l1ii_dataout;
	assign		wire_ni0ilOi_dataout = (n0OOO1i === 1'b1) ? wire_ni1l1lO_dataout : wire_ni0l1il_dataout;
	assign		wire_ni0ilOl_dataout = (n0OOO1i === 1'b1) ? wire_ni1l1Oi_dataout : wire_ni0l1iO_dataout;
	assign		wire_ni0ilOO_dataout = (n0OOO1i === 1'b1) ? wire_ni1l1Ol_dataout : wire_ni0l1li_dataout;
	assign		wire_ni0iO0i_dataout = (n0OOO1i === 1'b1) ? wire_ni1l01O_dataout : wire_ni0l1Ol_dataout;
	assign		wire_ni0iO0l_dataout = (n0OOO1i === 1'b1) ? wire_ni1l00i_dataout : wire_ni0l1OO_dataout;
	assign		wire_ni0iO0O_dataout = (n0OOO1i === 1'b1) ? wire_ni1l00l_dataout : wire_ni0l01i_dataout;
	assign		wire_ni0iO1i_dataout = (n0OOO1i === 1'b1) ? wire_ni1l1OO_dataout : wire_ni0l1ll_dataout;
	assign		wire_ni0iO1l_dataout = (n0OOO1i === 1'b1) ? wire_ni1l01i_dataout : wire_ni0l1lO_dataout;
	assign		wire_ni0iO1O_dataout = (n0OOO1i === 1'b1) ? wire_ni1l01l_dataout : wire_ni0l1Oi_dataout;
	assign		wire_ni0iOii_dataout = (n0OOO1i === 1'b1) ? wire_ni1l00O_dataout : wire_ni0l01l_dataout;
	assign		wire_ni0iOil_dataout = (n0OOO1i === 1'b1) ? wire_ni1l0ii_dataout : wire_ni0l01O_dataout;
	assign		wire_ni0iOiO_dataout = (n0OOO1i === 1'b1) ? wire_ni1l0il_dataout : wire_ni0l00i_dataout;
	assign		wire_ni0iOli_dataout = (n0OOO1i === 1'b1) ? wire_ni1l0iO_dataout : wire_ni0l00l_dataout;
	assign		wire_ni0iOll_dataout = (n0OOO1i === 1'b1) ? wire_ni1l0li_dataout : wire_ni0l00O_dataout;
	assign		wire_ni0iOlO_dataout = (n0OOO1i === 1'b1) ? wire_ni1l0ll_dataout : wire_ni0l0ii_dataout;
	assign		wire_ni0iOOi_dataout = (n0OOO1i === 1'b1) ? wire_ni1l0lO_dataout : wire_ni0l0il_dataout;
	assign		wire_ni0iOOl_dataout = (n0OOO0l === 1'b1) ? ni00iOl : ni0000i;
	assign		wire_ni0iOOO_dataout = (n0OOO0l === 1'b1) ? ni00iOO : ni0000l;
	assign		wire_ni0l00i_dataout = (n0OOO0l === 1'b1) ? ni00O0i : ni00iiO;
	assign		wire_ni0l00l_dataout = (n0OOO0l === 1'b1) ? ni00O0l : ni00ili;
	assign		wire_ni0l00O_dataout = (n0OOO0l === 1'b1) ? ni00O0O : ni00ill;
	assign		wire_ni0l01i_dataout = (n0OOO0l === 1'b1) ? ni00O1i : ni00i0O;
	assign		wire_ni0l01l_dataout = (n0OOO0l === 1'b1) ? ni00O1l : ni00iii;
	assign		wire_ni0l01O_dataout = (n0OOO0l === 1'b1) ? ni00O1O : ni00iil;
	assign		wire_ni0l0ii_dataout = (n0OOO0l === 1'b1) ? ni00Oii : ni00ilO;
	assign		wire_ni0l0il_dataout = (n0OOO0l === 1'b1) ? ni00Oil : ni00iOi;
	assign		wire_ni0l0Oi_dataout = (n0OOO1O === 1'b1) ? wire_ni1l11O_dataout : wire_ni0llil_dataout;
	assign		wire_ni0l0Ol_dataout = (n0OOO1O === 1'b1) ? wire_ni1l10i_dataout : wire_ni0lliO_dataout;
	assign		wire_ni0l0OO_dataout = (n0OOO1O === 1'b1) ? wire_ni1l10l_dataout : wire_ni0llli_dataout;
	assign		wire_ni0l10i_dataout = (n0OOO0l === 1'b1) ? ni00l0i : ni000iO;
	assign		wire_ni0l10l_dataout = (n0OOO0l === 1'b1) ? ni00l0l : ni000li;
	assign		wire_ni0l10O_dataout = (n0OOO0l === 1'b1) ? ni00l0O : ni000ll;
	assign		wire_ni0l11i_dataout = (n0OOO0l === 1'b1) ? ni00l1i : ni0000O;
	assign		wire_ni0l11l_dataout = (n0OOO0l === 1'b1) ? ni00l1l : ni000ii;
	assign		wire_ni0l11O_dataout = (n0OOO0l === 1'b1) ? ni00l1O : ni000il;
	assign		wire_ni0l1ii_dataout = (n0OOO0l === 1'b1) ? ni00lii : ni000lO;
	assign		wire_ni0l1il_dataout = (n0OOO0l === 1'b1) ? ni00lil : ni000Oi;
	assign		wire_ni0l1iO_dataout = (n0OOO0l === 1'b1) ? ni00liO : ni000Ol;
	assign		wire_ni0l1li_dataout = (n0OOO0l === 1'b1) ? ni00lli : ni000OO;
	assign		wire_ni0l1ll_dataout = (n0OOO0l === 1'b1) ? ni00lll : ni00i1i;
	assign		wire_ni0l1lO_dataout = (n0OOO0l === 1'b1) ? ni00llO : ni00i1l;
	assign		wire_ni0l1Oi_dataout = (n0OOO0l === 1'b1) ? ni00lOi : ni00i1O;
	assign		wire_ni0l1Ol_dataout = (n0OOO0l === 1'b1) ? ni00lOl : ni00i0i;
	assign		wire_ni0l1OO_dataout = (n0OOO0l === 1'b1) ? ni00lOO : ni00i0l;
	assign		wire_ni0li0i_dataout = (n0OOO1O === 1'b1) ? wire_ni1l1iO_dataout : wire_ni0llOl_dataout;
	assign		wire_ni0li0l_dataout = (n0OOO1O === 1'b1) ? wire_ni1l1li_dataout : wire_ni0llOO_dataout;
	assign		wire_ni0li0O_dataout = (n0OOO1O === 1'b1) ? wire_ni1l1ll_dataout : wire_ni0lO1i_dataout;
	assign		wire_ni0li1i_dataout = (n0OOO1O === 1'b1) ? wire_ni1l10O_dataout : wire_ni0llll_dataout;
	assign		wire_ni0li1l_dataout = (n0OOO1O === 1'b1) ? wire_ni1l1ii_dataout : wire_ni0lllO_dataout;
	assign		wire_ni0li1O_dataout = (n0OOO1O === 1'b1) ? wire_ni1l1il_dataout : wire_ni0llOi_dataout;
	assign		wire_ni0liii_dataout = (n0OOO1O === 1'b1) ? wire_ni1l1lO_dataout : wire_ni0lO1l_dataout;
	assign		wire_ni0liil_dataout = (n0OOO1O === 1'b1) ? wire_ni1l1Oi_dataout : wire_ni0lO1O_dataout;
	assign		wire_ni0liiO_dataout = (n0OOO1O === 1'b1) ? wire_ni1l1Ol_dataout : wire_ni0lO0i_dataout;
	assign		wire_ni0lili_dataout = (n0OOO1O === 1'b1) ? wire_ni1l1OO_dataout : wire_ni0lO0l_dataout;
	assign		wire_ni0lill_dataout = (n0OOO1O === 1'b1) ? wire_ni1l01i_dataout : wire_ni0lO0O_dataout;
	assign		wire_ni0lilO_dataout = (n0OOO1O === 1'b1) ? wire_ni1l01l_dataout : wire_ni0lOii_dataout;
	assign		wire_ni0liOi_dataout = (n0OOO1O === 1'b1) ? wire_ni1l01O_dataout : wire_ni0lOil_dataout;
	assign		wire_ni0liOl_dataout = (n0OOO1O === 1'b1) ? wire_ni1l00i_dataout : wire_ni0lOiO_dataout;
	assign		wire_ni0liOO_dataout = (n0OOO1O === 1'b1) ? wire_ni1l00l_dataout : wire_ni0lOli_dataout;
	assign		wire_ni0ll0i_dataout = (n0OOO1O === 1'b1) ? wire_ni1l0iO_dataout : wire_ni0lOOl_dataout;
	assign		wire_ni0ll0l_dataout = (n0OOO1O === 1'b1) ? wire_ni1l0li_dataout : wire_ni0lOOO_dataout;
	assign		wire_ni0ll0O_dataout = (n0OOO1O === 1'b1) ? wire_ni1l0ll_dataout : wire_ni0O11i_dataout;
	assign		wire_ni0ll1i_dataout = (n0OOO1O === 1'b1) ? wire_ni1l00O_dataout : wire_ni0lOll_dataout;
	assign		wire_ni0ll1l_dataout = (n0OOO1O === 1'b1) ? wire_ni1l0ii_dataout : wire_ni0lOlO_dataout;
	assign		wire_ni0ll1O_dataout = (n0OOO1O === 1'b1) ? wire_ni1l0il_dataout : wire_ni0lOOi_dataout;
	assign		wire_ni0llii_dataout = (n0OOO1O === 1'b1) ? wire_ni1l0lO_dataout : wire_ni0O11l_dataout;
	assign		wire_ni0llil_dataout = (n0OOO0l === 1'b1) ? ni0000i : ni0il1O;
	assign		wire_ni0lliO_dataout = (n0OOO0l === 1'b1) ? ni0000l : ni01Oli;
	assign		wire_ni0llli_dataout = (n0OOO0l === 1'b1) ? ni0000O : ni01Oll;
	assign		wire_ni0llll_dataout = (n0OOO0l === 1'b1) ? ni000ii : ni01OlO;
	assign		wire_ni0lllO_dataout = (n0OOO0l === 1'b1) ? ni000il : ni01OOi;
	assign		wire_ni0llOi_dataout = (n0OOO0l === 1'b1) ? ni000iO : ni01OOl;
	assign		wire_ni0llOl_dataout = (n0OOO0l === 1'b1) ? ni000li : ni01OOO;
	assign		wire_ni0llOO_dataout = (n0OOO0l === 1'b1) ? ni000ll : ni0011i;
	assign		wire_ni0lO0i_dataout = (n0OOO0l === 1'b1) ? ni000OO : ni0010l;
	assign		wire_ni0lO0l_dataout = (n0OOO0l === 1'b1) ? ni00i1i : ni0010O;
	assign		wire_ni0lO0O_dataout = (n0OOO0l === 1'b1) ? ni00i1l : ni001ii;
	assign		wire_ni0lO1i_dataout = (n0OOO0l === 1'b1) ? ni000lO : ni0011l;
	assign		wire_ni0lO1l_dataout = (n0OOO0l === 1'b1) ? ni000Oi : ni0011O;
	assign		wire_ni0lO1O_dataout = (n0OOO0l === 1'b1) ? ni000Ol : ni0010i;
	assign		wire_ni0lOii_dataout = (n0OOO0l === 1'b1) ? ni00i1O : ni001il;
	assign		wire_ni0lOil_dataout = (n0OOO0l === 1'b1) ? ni00i0i : ni001iO;
	assign		wire_ni0lOiO_dataout = (n0OOO0l === 1'b1) ? ni00i0l : ni001li;
	assign		wire_ni0lOli_dataout = (n0OOO0l === 1'b1) ? ni00i0O : ni001ll;
	assign		wire_ni0lOll_dataout = (n0OOO0l === 1'b1) ? ni00iii : ni001lO;
	assign		wire_ni0lOlO_dataout = (n0OOO0l === 1'b1) ? ni00iil : ni001Oi;
	assign		wire_ni0lOOi_dataout = (n0OOO0l === 1'b1) ? ni00iiO : ni001Ol;
	assign		wire_ni0lOOl_dataout = (n0OOO0l === 1'b1) ? ni00ili : ni001OO;
	assign		wire_ni0lOOO_dataout = (n0OOO0l === 1'b1) ? ni00ill : ni0001i;
	assign		wire_ni0O11i_dataout = (n0OOO0l === 1'b1) ? ni00ilO : ni0001l;
	assign		wire_ni0O11l_dataout = (n0OOO0l === 1'b1) ? ni00iOi : ni0001O;
	assign		wire_ni0O1il_dataout = ((~ n0OOOil) === 1'b1) ? n0OOOii : ni0Oi0i;
	assign		wire_ni0Oi0O_dataout = (((~ n0OOOiO) & n0OOOii) === 1'b1) ? wire_ni0Oili_o[1] : wire_ni0Oiii_dataout;
	assign		wire_ni0Oiii_dataout = ((n0OOOiO & (~ n0OOOii)) === 1'b1) ? wire_ni0Oiil_o[0] : ni0Oi1O;
	assign		wire_ni0OilO_dataout = (ni0Oi0l === 1'b1) ? ni0il1O : nii110i;
	assign		wire_ni0OiOi_dataout = (ni0Oi0l === 1'b1) ? ni01Oli : ni0O1iO;
	assign		wire_ni0OiOl_dataout = (ni0Oi0l === 1'b1) ? ni01Oll : ni0O1li;
	assign		wire_ni0OiOO_dataout = (ni0Oi0l === 1'b1) ? ni01OlO : ni0O1ll;
	assign		wire_ni0Ol0i_dataout = (ni0Oi0l === 1'b1) ? ni0011i : ni0O1OO;
	assign		wire_ni0Ol0l_dataout = (ni0Oi0l === 1'b1) ? ni0011l : ni0O01i;
	assign		wire_ni0Ol0O_dataout = (ni0Oi0l === 1'b1) ? ni0011O : ni0O01l;
	assign		wire_ni0Ol1i_dataout = (ni0Oi0l === 1'b1) ? ni01OOi : ni0O1lO;
	assign		wire_ni0Ol1l_dataout = (ni0Oi0l === 1'b1) ? ni01OOl : ni0O1Oi;
	assign		wire_ni0Ol1O_dataout = (ni0Oi0l === 1'b1) ? ni01OOO : ni0O1Ol;
	assign		wire_ni0Olii_dataout = (ni0Oi0l === 1'b1) ? ni0010i : ni0O01O;
	assign		wire_ni0Olil_dataout = (ni0Oi0l === 1'b1) ? ni0010l : ni0O00i;
	assign		wire_ni0OliO_dataout = (ni0Oi0l === 1'b1) ? ni0010O : ni0O00l;
	assign		wire_ni0Olli_dataout = (ni0Oi0l === 1'b1) ? ni001ii : ni0O00O;
	assign		wire_ni0Olll_dataout = (ni0Oi0l === 1'b1) ? ni001il : ni0O0ii;
	assign		wire_ni0OllO_dataout = (ni0Oi0l === 1'b1) ? ni001iO : ni0O0il;
	assign		wire_ni0OlOi_dataout = (ni0Oi0l === 1'b1) ? ni001li : ni0O0iO;
	assign		wire_ni0OlOl_dataout = (ni0Oi0l === 1'b1) ? ni001ll : ni0O0li;
	assign		wire_ni0OlOO_dataout = (ni0Oi0l === 1'b1) ? ni001lO : ni0O0ll;
	assign		wire_ni0OO0i_dataout = (ni0Oi0l === 1'b1) ? ni0001i : ni0O0OO;
	assign		wire_ni0OO0l_dataout = (ni0Oi0l === 1'b1) ? ni0001l : ni0Oi1i;
	assign		wire_ni0OO0O_dataout = (ni0Oi0l === 1'b1) ? ni0001O : ni0Oi1l;
	assign		wire_ni0OO1i_dataout = (ni0Oi0l === 1'b1) ? ni001Oi : ni0O0lO;
	assign		wire_ni0OO1l_dataout = (ni0Oi0l === 1'b1) ? ni001Ol : ni0O0Oi;
	assign		wire_ni0OO1O_dataout = (ni0Oi0l === 1'b1) ? ni001OO : ni0O0Ol;
	assign		wire_ni1l00i_dataout = (n0OOili === 1'b1) ? nl11i1O : wire_ni1liOl_dataout;
	assign		wire_ni1l00l_dataout = (n0OOili === 1'b1) ? nl11i0i : wire_ni1liOO_dataout;
	assign		wire_ni1l00O_dataout = (n0OOili === 1'b1) ? nl11i0l : wire_ni1ll1i_dataout;
	assign		wire_ni1l01i_dataout = (n0OOili === 1'b1) ? nl110OO : wire_ni1lill_dataout;
	assign		wire_ni1l01l_dataout = (n0OOili === 1'b1) ? nl11i1i : wire_ni1lilO_dataout;
	assign		wire_ni1l01O_dataout = (n0OOili === 1'b1) ? nl11i1l : wire_ni1liOi_dataout;
	assign		wire_ni1l0ii_dataout = (n0OOili === 1'b1) ? nl11i0O : wire_ni1ll1l_dataout;
	assign		wire_ni1l0il_dataout = (n0OOili === 1'b1) ? nl11iii : wire_ni1ll1O_dataout;
	assign		wire_ni1l0iO_dataout = (n0OOili === 1'b1) ? nl11iil : wire_ni1ll0i_dataout;
	assign		wire_ni1l0li_dataout = (n0OOili === 1'b1) ? nl11iiO : wire_ni1ll0l_dataout;
	assign		wire_ni1l0ll_dataout = (n0OOili === 1'b1) ? nl11ill : wire_ni1ll0O_dataout;
	assign		wire_ni1l0lO_dataout = (n0OOili === 1'b1) ? nli11lO : wire_ni1llii_dataout;
	and(wire_ni1l0Oi_dataout, wire_ni1llil_dataout, ~(n0OOill));
	and(wire_ni1l0Ol_dataout, wire_ni1lliO_dataout, ~(n0OOill));
	and(wire_ni1l0OO_dataout, wire_ni1llli_dataout, ~(n0OOill));
	assign		wire_ni1l10i_dataout = (n0OOili === 1'b1) ? nl1101O : wire_ni1l0Ol_dataout;
	assign		wire_ni1l10l_dataout = (n0OOili === 1'b1) ? nl1100i : wire_ni1l0OO_dataout;
	assign		wire_ni1l10O_dataout = (n0OOili === 1'b1) ? nl1100l : wire_ni1li1i_dataout;
	assign		wire_ni1l11O_dataout = (n0OOili === 1'b1) ? nl1101l : wire_ni1l0Oi_dataout;
	assign		wire_ni1l1ii_dataout = (n0OOili === 1'b1) ? nl1100O : wire_ni1li1l_dataout;
	assign		wire_ni1l1il_dataout = (n0OOili === 1'b1) ? nl110ii : wire_ni1li1O_dataout;
	assign		wire_ni1l1iO_dataout = (n0OOili === 1'b1) ? nl110il : wire_ni1li0i_dataout;
	assign		wire_ni1l1li_dataout = (n0OOili === 1'b1) ? nl110iO : wire_ni1li0l_dataout;
	assign		wire_ni1l1ll_dataout = (n0OOili === 1'b1) ? nl110li : wire_ni1li0O_dataout;
	assign		wire_ni1l1lO_dataout = (n0OOili === 1'b1) ? nl110ll : wire_ni1liii_dataout;
	assign		wire_ni1l1Oi_dataout = (n0OOili === 1'b1) ? nl110lO : wire_ni1liil_dataout;
	assign		wire_ni1l1Ol_dataout = (n0OOili === 1'b1) ? nl110Oi : wire_ni1liiO_dataout;
	assign		wire_ni1l1OO_dataout = (n0OOili === 1'b1) ? nl110Ol : wire_ni1lili_dataout;
	and(wire_ni1li0i_dataout, wire_ni1llOl_dataout, ~(n0OOill));
	and(wire_ni1li0l_dataout, wire_ni1llOO_dataout, ~(n0OOill));
	and(wire_ni1li0O_dataout, wire_ni1lO1i_dataout, ~(n0OOill));
	and(wire_ni1li1i_dataout, wire_ni1llll_dataout, ~(n0OOill));
	and(wire_ni1li1l_dataout, wire_ni1lllO_dataout, ~(n0OOill));
	and(wire_ni1li1O_dataout, wire_ni1llOi_dataout, ~(n0OOill));
	and(wire_ni1liii_dataout, wire_ni1lO1l_dataout, ~(n0OOill));
	and(wire_ni1liil_dataout, wire_ni1lO1O_dataout, ~(n0OOill));
	and(wire_ni1liiO_dataout, wire_ni1lO0i_dataout, ~(n0OOill));
	and(wire_ni1lili_dataout, wire_ni1lO0l_dataout, ~(n0OOill));
	and(wire_ni1lill_dataout, wire_ni1lO0O_dataout, ~(n0OOill));
	and(wire_ni1lilO_dataout, wire_ni1lOii_dataout, ~(n0OOill));
	and(wire_ni1liOi_dataout, wire_ni1lOil_dataout, ~(n0OOill));
	and(wire_ni1liOl_dataout, wire_ni1lOiO_dataout, ~(n0OOill));
	and(wire_ni1liOO_dataout, wire_ni1lOli_dataout, ~(n0OOill));
	and(wire_ni1ll0i_dataout, wire_ni1lOOl_dataout, ~(n0OOill));
	and(wire_ni1ll0l_dataout, wire_ni1lOOO_dataout, ~(n0OOill));
	and(wire_ni1ll0O_dataout, wire_ni1O11i_dataout, ~(n0OOill));
	and(wire_ni1ll1i_dataout, wire_ni1lOll_dataout, ~(n0OOill));
	and(wire_ni1ll1l_dataout, wire_ni1lOlO_dataout, ~(n0OOill));
	and(wire_ni1ll1O_dataout, wire_ni1lOOi_dataout, ~(n0OOill));
	assign		wire_ni1llii_dataout = (n0OOill === 1'b1) ? nii00li : wire_ni1O11l_dataout;
	assign		wire_ni1llil_dataout = (n0OOilO === 1'b1) ? nl1iO1l : wire_ni1O11O_dataout;
	assign		wire_ni1lliO_dataout = (n0OOilO === 1'b1) ? nl1iO1O : wire_ni1O10i_dataout;
	assign		wire_ni1llli_dataout = (n0OOilO === 1'b1) ? nl1iO0i : wire_ni1O10l_dataout;
	assign		wire_ni1llll_dataout = (n0OOilO === 1'b1) ? nl1iO0l : wire_ni1O10O_dataout;
	assign		wire_ni1lllO_dataout = (n0OOilO === 1'b1) ? nl1iO0O : wire_ni1O1ii_dataout;
	assign		wire_ni1llOi_dataout = (n0OOilO === 1'b1) ? nl1iOii : wire_ni1O1il_dataout;
	assign		wire_ni1llOl_dataout = (n0OOilO === 1'b1) ? nl1iOil : wire_ni1O1iO_dataout;
	assign		wire_ni1llOO_dataout = (n0OOilO === 1'b1) ? nl1iOli : wire_ni1O1li_dataout;
	assign		wire_ni1lO0i_dataout = (n0OOilO === 1'b1) ? nl1l11i : wire_ni1O1Ol_dataout;
	assign		wire_ni1lO0l_dataout = (n0OOilO === 1'b1) ? nl1l11l : wire_ni1O1OO_dataout;
	assign		wire_ni1lO0O_dataout = (n0OOilO === 1'b1) ? nl1l11O : wire_ni1O01i_dataout;
	assign		wire_ni1lO1i_dataout = (n0OOilO === 1'b1) ? nl1iOOi : wire_ni1O1ll_dataout;
	assign		wire_ni1lO1l_dataout = (n0OOilO === 1'b1) ? nl1iOOl : wire_ni1O1lO_dataout;
	assign		wire_ni1lO1O_dataout = (n0OOilO === 1'b1) ? nl1iOOO : wire_ni1O1Oi_dataout;
	assign		wire_ni1lOii_dataout = (n0OOilO === 1'b1) ? nl1l10i : wire_ni1O01l_dataout;
	assign		wire_ni1lOil_dataout = (n0OOilO === 1'b1) ? nl1l10O : wire_ni1O01O_dataout;
	assign		wire_ni1lOiO_dataout = (n0OOilO === 1'b1) ? nl1l1iO : wire_ni1O00i_dataout;
	assign		wire_ni1lOli_dataout = (n0OOilO === 1'b1) ? nl1l1li : wire_ni1O00l_dataout;
	assign		wire_ni1lOll_dataout = (n0OOilO === 1'b1) ? nl1l1ll : wire_ni1O00O_dataout;
	assign		wire_ni1lOlO_dataout = (n0OOilO === 1'b1) ? nl1l1lO : wire_ni1O0ii_dataout;
	assign		wire_ni1lOOi_dataout = (n0OOilO === 1'b1) ? nl1l1Oi : wire_ni1O0il_dataout;
	assign		wire_ni1lOOl_dataout = (n0OOilO === 1'b1) ? nl1l1Ol : wire_ni1O0iO_dataout;
	assign		wire_ni1lOOO_dataout = (n0OOilO === 1'b1) ? nl1l1OO : wire_ni1O0li_dataout;
	assign		wire_ni1O00i_dataout = (n0OOiOi === 1'b1) ? nl11i1O : wire_ni1OiOl_dataout;
	assign		wire_ni1O00l_dataout = (n0OOiOi === 1'b1) ? nl11i0i : wire_ni1OiOO_dataout;
	assign		wire_ni1O00O_dataout = (n0OOiOi === 1'b1) ? nl11i0l : wire_ni1Ol1i_dataout;
	assign		wire_ni1O01i_dataout = (n0OOiOi === 1'b1) ? nl110OO : wire_ni1Oill_dataout;
	assign		wire_ni1O01l_dataout = (n0OOiOi === 1'b1) ? nl11i1i : wire_ni1OilO_dataout;
	assign		wire_ni1O01O_dataout = (n0OOiOi === 1'b1) ? nl11i1l : wire_ni1OiOi_dataout;
	assign		wire_ni1O0ii_dataout = (n0OOiOi === 1'b1) ? nl11i0O : wire_ni1Ol1l_dataout;
	assign		wire_ni1O0il_dataout = (n0OOiOi === 1'b1) ? nl11iii : wire_ni1Ol1O_dataout;
	assign		wire_ni1O0iO_dataout = (n0OOiOi === 1'b1) ? nl11iil : wire_ni1Ol0i_dataout;
	assign		wire_ni1O0li_dataout = (n0OOiOi === 1'b1) ? nl11iiO : wire_ni1Ol0l_dataout;
	assign		wire_ni1O0ll_dataout = (n0OOiOi === 1'b1) ? nl11ill : wire_ni1Ol0O_dataout;
	assign		wire_ni1O0lO_dataout = (n0OOiOi === 1'b1) ? nii00li : wire_ni1Olii_dataout;
	assign		wire_ni1O0Oi_dataout = (n0OOiOl === 1'b1) ? nl100iO : wire_ni1Olil_dataout;
	assign		wire_ni1O0Ol_dataout = (n0OOiOl === 1'b1) ? nl100li : wire_ni1OliO_dataout;
	assign		wire_ni1O0OO_dataout = (n0OOiOl === 1'b1) ? nl100ll : wire_ni1Olli_dataout;
	assign		wire_ni1O10i_dataout = (n0OOiOi === 1'b1) ? nl1101O : wire_ni1O0Ol_dataout;
	assign		wire_ni1O10l_dataout = (n0OOiOi === 1'b1) ? nl1100i : wire_ni1O0OO_dataout;
	assign		wire_ni1O10O_dataout = (n0OOiOi === 1'b1) ? nl1100l : wire_ni1Oi1i_dataout;
	assign		wire_ni1O11i_dataout = (n0OOilO === 1'b1) ? nl1l01l : wire_ni1O0ll_dataout;
	assign		wire_ni1O11l_dataout = (n0OOilO === 1'b1) ? nli1ilO : wire_ni1O0lO_dataout;
	assign		wire_ni1O11O_dataout = (n0OOiOi === 1'b1) ? nl1101l : wire_ni1O0Oi_dataout;
	assign		wire_ni1O1ii_dataout = (n0OOiOi === 1'b1) ? nl1100O : wire_ni1Oi1l_dataout;
	assign		wire_ni1O1il_dataout = (n0OOiOi === 1'b1) ? nl110ii : wire_ni1Oi1O_dataout;
	assign		wire_ni1O1iO_dataout = (n0OOiOi === 1'b1) ? nl110il : wire_ni1Oi0i_dataout;
	assign		wire_ni1O1li_dataout = (n0OOiOi === 1'b1) ? nl110iO : wire_ni1Oi0l_dataout;
	assign		wire_ni1O1ll_dataout = (n0OOiOi === 1'b1) ? nl110li : wire_ni1Oi0O_dataout;
	assign		wire_ni1O1lO_dataout = (n0OOiOi === 1'b1) ? nl110ll : wire_ni1Oiii_dataout;
	assign		wire_ni1O1Oi_dataout = (n0OOiOi === 1'b1) ? nl110lO : wire_ni1Oiil_dataout;
	assign		wire_ni1O1Ol_dataout = (n0OOiOi === 1'b1) ? nl110Oi : wire_ni1OiiO_dataout;
	assign		wire_ni1O1OO_dataout = (n0OOiOi === 1'b1) ? nl110Ol : wire_ni1Oili_dataout;
	assign		wire_ni1Oi0i_dataout = (n0OOiOl === 1'b1) ? nl100OO : wire_ni1OlOl_dataout;
	assign		wire_ni1Oi0l_dataout = (n0OOiOl === 1'b1) ? nl10i1i : wire_ni1OlOO_dataout;
	assign		wire_ni1Oi0O_dataout = (n0OOiOl === 1'b1) ? nl10i1l : wire_ni1OO1i_dataout;
	assign		wire_ni1Oi1i_dataout = (n0OOiOl === 1'b1) ? nl100lO : wire_ni1Olll_dataout;
	assign		wire_ni1Oi1l_dataout = (n0OOiOl === 1'b1) ? nl100Oi : wire_ni1OllO_dataout;
	assign		wire_ni1Oi1O_dataout = (n0OOiOl === 1'b1) ? nl100Ol : wire_ni1OlOi_dataout;
	assign		wire_ni1Oiii_dataout = (n0OOiOl === 1'b1) ? nl10i1O : wire_ni1OO1l_dataout;
	assign		wire_ni1Oiil_dataout = (n0OOiOl === 1'b1) ? nl10i0i : wire_ni1OO1O_dataout;
	assign		wire_ni1OiiO_dataout = (n0OOiOl === 1'b1) ? nl10i0l : wire_ni1OO0i_dataout;
	assign		wire_ni1Oili_dataout = (n0OOiOl === 1'b1) ? nl10i0O : wire_ni1OO0l_dataout;
	assign		wire_ni1Oill_dataout = (n0OOiOl === 1'b1) ? nl10iii : wire_ni1OO0O_dataout;
	assign		wire_ni1OilO_dataout = (n0OOiOl === 1'b1) ? nl10iil : wire_ni1OOii_dataout;
	assign		wire_ni1OiOi_dataout = (n0OOiOl === 1'b1) ? nl10iiO : wire_ni1OOil_dataout;
	assign		wire_ni1OiOl_dataout = (n0OOiOl === 1'b1) ? nl10ili : wire_ni1OOiO_dataout;
	assign		wire_ni1OiOO_dataout = (n0OOiOl === 1'b1) ? nl10ill : wire_ni1OOli_dataout;
	assign		wire_ni1Ol0i_dataout = (n0OOiOl === 1'b1) ? nl10iOO : wire_ni1OOOl_dataout;
	assign		wire_ni1Ol0l_dataout = (n0OOiOl === 1'b1) ? nl10l1i : wire_ni1OOOO_dataout;
	assign		wire_ni1Ol0O_dataout = (n0OOiOl === 1'b1) ? nl10l1O : wire_ni0111i_dataout;
	assign		wire_ni1Ol1i_dataout = (n0OOiOl === 1'b1) ? nl10ilO : wire_ni1OOll_dataout;
	assign		wire_ni1Ol1l_dataout = (n0OOiOl === 1'b1) ? nl10iOi : wire_ni1OOlO_dataout;
	assign		wire_ni1Ol1O_dataout = (n0OOiOl === 1'b1) ? nl10iOl : wire_ni1OOOi_dataout;
	assign		wire_ni1Olii_dataout = (n0OOiOl === 1'b1) ? nil10lO : wire_ni0111l_dataout;
	and(wire_ni1Olil_dataout, nl100iO, n0OOiOO);
	and(wire_ni1OliO_dataout, nl100li, n0OOiOO);
	and(wire_ni1Olli_dataout, nl100ll, n0OOiOO);
	and(wire_ni1Olll_dataout, nl100lO, n0OOiOO);
	and(wire_ni1OllO_dataout, nl100Oi, n0OOiOO);
	and(wire_ni1OlOi_dataout, nl100Ol, n0OOiOO);
	and(wire_ni1OlOl_dataout, nl100OO, n0OOiOO);
	and(wire_ni1OlOO_dataout, nl10i1i, n0OOiOO);
	and(wire_ni1OO0i_dataout, nl10i0l, n0OOiOO);
	and(wire_ni1OO0l_dataout, nl10i0O, n0OOiOO);
	and(wire_ni1OO0O_dataout, nl10iii, n0OOiOO);
	and(wire_ni1OO1i_dataout, nl10i1l, n0OOiOO);
	and(wire_ni1OO1l_dataout, nl10i1O, n0OOiOO);
	and(wire_ni1OO1O_dataout, nl10i0i, n0OOiOO);
	and(wire_ni1OOii_dataout, nl10iil, n0OOiOO);
	and(wire_ni1OOil_dataout, nl10iiO, n0OOiOO);
	and(wire_ni1OOiO_dataout, nl10ili, n0OOiOO);
	and(wire_ni1OOli_dataout, nl10ill, n0OOiOO);
	and(wire_ni1OOll_dataout, nl10ilO, n0OOiOO);
	and(wire_ni1OOlO_dataout, nl10iOi, n0OOiOO);
	and(wire_ni1OOOi_dataout, nl10iOl, n0OOiOO);
	and(wire_ni1OOOl_dataout, nl10iOO, n0OOiOO);
	and(wire_ni1OOOO_dataout, nl10l1i, n0OOiOO);
	and(wire_nii001i_dataout, wire_nii001l_o[6], ~(n00il));
	assign		wire_nii00ll_dataout = (nil101O === 1'b1) ? wire_nii00Ol_dataout : wire_nii00lO_dataout;
	or(wire_nii00lO_dataout, wire_nii00Oi_dataout, ni111Ol);
	assign		wire_nii00Oi_dataout = (ni111Oi === 1'b1) ? (~ nii0lOi) : (~ nii0lOl);
	assign		wire_nii00Ol_dataout = (ni111Ol === 1'b1) ? (~ nii0lOl) : wire_nii00OO_dataout;
	assign		wire_nii00OO_dataout = (ni111Oi === 1'b1) ? (~ nii0lll) : (~ nii0lOi);
	and(wire_nii011i_dataout, wire_nii011l_o[4], ~(wire_nii1O0O_o));
	or(wire_nii01ll_dataout, wire_nii001l_o[1], n00il);
	and(wire_nii01lO_dataout, wire_nii001l_o[2], ~(n00il));
	and(wire_nii01Oi_dataout, wire_nii001l_o[3], ~(n00il));
	and(wire_nii01Ol_dataout, wire_nii001l_o[4], ~(n00il));
	and(wire_nii01OO_dataout, wire_nii001l_o[5], ~(n00il));
	and(wire_nii1OOi_dataout, wire_nii011l_o[1], ~(wire_nii1O0O_o));
	and(wire_nii1OOl_dataout, wire_nii011l_o[2], ~(wire_nii1O0O_o));
	and(wire_nii1OOO_dataout, wire_nii011l_o[3], ~(wire_nii1O0O_o));
	assign		wire_niiiO0i_dataout = (ni111il === 1'b1) ? din_0_data[1] : wire_niil1Ol_dataout;
	assign		wire_niiiO0l_dataout = (ni111il === 1'b1) ? din_0_data[2] : wire_niil1OO_dataout;
	assign		wire_niiiO0O_dataout = (ni111il === 1'b1) ? din_0_data[3] : wire_niil01i_dataout;
	or(wire_niiiO1i_dataout, wire_niiiO1l_dataout, ni111il);
	and(wire_niiiO1l_dataout, nii0lOl, ~(ni111OO));
	assign		wire_niiiO1O_dataout = (ni111il === 1'b1) ? din_0_data[0] : wire_niil1Oi_dataout;
	assign		wire_niiiOii_dataout = (ni111il === 1'b1) ? din_0_data[4] : wire_niil01l_dataout;
	assign		wire_niiiOil_dataout = (ni111il === 1'b1) ? din_0_data[5] : wire_niil01O_dataout;
	assign		wire_niiiOiO_dataout = (ni111il === 1'b1) ? din_0_data[6] : wire_niil00i_dataout;
	assign		wire_niiiOli_dataout = (ni111il === 1'b1) ? din_0_data[7] : wire_niil00l_dataout;
	assign		wire_niiiOll_dataout = (ni111il === 1'b1) ? din_0_data[8] : wire_niil00O_dataout;
	assign		wire_niiiOlO_dataout = (ni111il === 1'b1) ? din_0_data[9] : wire_niil0ii_dataout;
	assign		wire_niiiOOi_dataout = (ni111il === 1'b1) ? din_0_data[10] : wire_niil0il_dataout;
	assign		wire_niiiOOl_dataout = (ni111il === 1'b1) ? din_0_data[11] : wire_niil0iO_dataout;
	assign		wire_niiiOOO_dataout = (ni111il === 1'b1) ? din_0_data[12] : wire_niil0li_dataout;
	or(wire_niil00i_dataout, niiiill, ni111OO);
	or(wire_niil00l_dataout, niiiilO, ni111OO);
	or(wire_niil00O_dataout, niiiiOi, ni111OO);
	or(wire_niil01i_dataout, niiiiil, ni111OO);
	or(wire_niil01l_dataout, niiiiiO, ni111OO);
	or(wire_niil01O_dataout, niiiili, ni111OO);
	or(wire_niil0ii_dataout, niiiiOl, ni111OO);
	or(wire_niil0il_dataout, niiiiOO, ni111OO);
	or(wire_niil0iO_dataout, niiil1i, ni111OO);
	or(wire_niil0li_dataout, niiil1l, ni111OO);
	or(wire_niil0ll_dataout, niiil1O, ni111OO);
	or(wire_niil0lO_dataout, niiil0i, ni111OO);
	or(wire_niil0Oi_dataout, niiil0l, ni111OO);
	or(wire_niil0Ol_dataout, niiil0O, ni111OO);
	or(wire_niil0OO_dataout, niiilii, ni111OO);
	assign		wire_niil10i_dataout = (ni111il === 1'b1) ? din_0_data[16] : wire_niil0Ol_dataout;
	assign		wire_niil10l_dataout = (ni111il === 1'b1) ? din_0_data[17] : wire_niil0OO_dataout;
	assign		wire_niil10O_dataout = (ni111il === 1'b1) ? din_0_data[18] : wire_niili1i_dataout;
	assign		wire_niil11i_dataout = (ni111il === 1'b1) ? din_0_data[13] : wire_niil0ll_dataout;
	assign		wire_niil11l_dataout = (ni111il === 1'b1) ? din_0_data[14] : wire_niil0lO_dataout;
	assign		wire_niil11O_dataout = (ni111il === 1'b1) ? din_0_data[15] : wire_niil0Oi_dataout;
	assign		wire_niil1ii_dataout = (ni111il === 1'b1) ? din_0_data[19] : wire_niili1l_dataout;
	assign		wire_niil1il_dataout = (ni111il === 1'b1) ? din_0_data[20] : wire_niili1O_dataout;
	assign		wire_niil1iO_dataout = (ni111il === 1'b1) ? din_0_data[21] : wire_niili0i_dataout;
	assign		wire_niil1li_dataout = (ni111il === 1'b1) ? din_0_data[22] : wire_niili0l_dataout;
	assign		wire_niil1ll_dataout = (ni111il === 1'b1) ? din_0_data[23] : wire_niili0O_dataout;
	assign		wire_niil1lO_dataout = (ni111il === 1'b1) ? din_0_endofpacket : wire_niiliii_dataout;
	or(wire_niil1Oi_dataout, niiii0l, ni111OO);
	or(wire_niil1Ol_dataout, niiii0O, ni111OO);
	or(wire_niil1OO_dataout, niiiiii, ni111OO);
	or(wire_niili0i_dataout, niiilll, ni111OO);
	or(wire_niili0l_dataout, niiillO, ni111OO);
	or(wire_niili0O_dataout, niiilOi, ni111OO);
	or(wire_niili1i_dataout, niiilil, ni111OO);
	or(wire_niili1l_dataout, niiiliO, ni111OO);
	or(wire_niili1O_dataout, niiilli, ni111OO);
	or(wire_niiliii_dataout, niiilOl, ni111OO);
	or(wire_niiliOi_dataout, wire_niiliOl_dataout, ni111iO);
	assign		wire_niiliOl_dataout = (ni111OO === 1'b1) ? nii0lOl : nii0lOi;
	assign		wire_niiliOO_dataout = (ni111iO === 1'b1) ? din_0_data[0] : wire_niilOli_dataout;
	assign		wire_niill0i_dataout = (ni111iO === 1'b1) ? din_0_data[4] : wire_niilOOl_dataout;
	assign		wire_niill0l_dataout = (ni111iO === 1'b1) ? din_0_data[5] : wire_niilOOO_dataout;
	assign		wire_niill0O_dataout = (ni111iO === 1'b1) ? din_0_data[6] : wire_niiO11i_dataout;
	assign		wire_niill1i_dataout = (ni111iO === 1'b1) ? din_0_data[1] : wire_niilOll_dataout;
	assign		wire_niill1l_dataout = (ni111iO === 1'b1) ? din_0_data[2] : wire_niilOlO_dataout;
	assign		wire_niill1O_dataout = (ni111iO === 1'b1) ? din_0_data[3] : wire_niilOOi_dataout;
	assign		wire_niillii_dataout = (ni111iO === 1'b1) ? din_0_data[7] : wire_niiO11l_dataout;
	assign		wire_niillil_dataout = (ni111iO === 1'b1) ? din_0_data[8] : wire_niiO11O_dataout;
	assign		wire_niilliO_dataout = (ni111iO === 1'b1) ? din_0_data[9] : wire_niiO10i_dataout;
	assign		wire_niillli_dataout = (ni111iO === 1'b1) ? din_0_data[10] : wire_niiO10l_dataout;
	assign		wire_niillll_dataout = (ni111iO === 1'b1) ? din_0_data[11] : wire_niiO10O_dataout;
	assign		wire_niilllO_dataout = (ni111iO === 1'b1) ? din_0_data[12] : wire_niiO1ii_dataout;
	assign		wire_niillOi_dataout = (ni111iO === 1'b1) ? din_0_data[13] : wire_niiO1il_dataout;
	assign		wire_niillOl_dataout = (ni111iO === 1'b1) ? din_0_data[14] : wire_niiO1iO_dataout;
	assign		wire_niillOO_dataout = (ni111iO === 1'b1) ? din_0_data[15] : wire_niiO1li_dataout;
	assign		wire_niilO0i_dataout = (ni111iO === 1'b1) ? din_0_data[19] : wire_niiO1Ol_dataout;
	assign		wire_niilO0l_dataout = (ni111iO === 1'b1) ? din_0_data[20] : wire_niiO1OO_dataout;
	assign		wire_niilO0O_dataout = (ni111iO === 1'b1) ? din_0_data[21] : wire_niiO01i_dataout;
	assign		wire_niilO1i_dataout = (ni111iO === 1'b1) ? din_0_data[16] : wire_niiO1ll_dataout;
	assign		wire_niilO1l_dataout = (ni111iO === 1'b1) ? din_0_data[17] : wire_niiO1lO_dataout;
	assign		wire_niilO1O_dataout = (ni111iO === 1'b1) ? din_0_data[18] : wire_niiO1Oi_dataout;
	assign		wire_niilOii_dataout = (ni111iO === 1'b1) ? din_0_data[22] : wire_niiO01l_dataout;
	assign		wire_niilOil_dataout = (ni111iO === 1'b1) ? din_0_data[23] : wire_niiO01O_dataout;
	assign		wire_niilOiO_dataout = (ni111iO === 1'b1) ? din_0_endofpacket : wire_niiO00i_dataout;
	assign		wire_niilOli_dataout = (ni111OO === 1'b1) ? niiii0l : niii1li;
	assign		wire_niilOll_dataout = (ni111OO === 1'b1) ? niiii0O : niii1ll;
	assign		wire_niilOlO_dataout = (ni111OO === 1'b1) ? niiiiii : niii1lO;
	assign		wire_niilOOi_dataout = (ni111OO === 1'b1) ? niiiiil : niii1Oi;
	assign		wire_niilOOl_dataout = (ni111OO === 1'b1) ? niiiiiO : niii1Ol;
	assign		wire_niilOOO_dataout = (ni111OO === 1'b1) ? niiiili : niii1OO;
	assign		wire_niiO00i_dataout = (ni111OO === 1'b1) ? niiilOl : niiii0i;
	assign		wire_niiO01i_dataout = (ni111OO === 1'b1) ? niiilll : niiii1i;
	assign		wire_niiO01l_dataout = (ni111OO === 1'b1) ? niiillO : niiii1l;
	assign		wire_niiO01O_dataout = (ni111OO === 1'b1) ? niiilOi : niiii1O;
	or(wire_niiO0iO_dataout, wire_niiO0li_dataout, ni111ll);
	assign		wire_niiO0li_dataout = (ni111OO === 1'b1) ? nii0lOi : nii0lll;
	assign		wire_niiO0ll_dataout = (ni111ll === 1'b1) ? din_0_data[0] : wire_niiOl0O_dataout;
	assign		wire_niiO0lO_dataout = (ni111ll === 1'b1) ? din_0_data[1] : wire_niiOlii_dataout;
	assign		wire_niiO0Oi_dataout = (ni111ll === 1'b1) ? din_0_data[2] : wire_niiOlil_dataout;
	assign		wire_niiO0Ol_dataout = (ni111ll === 1'b1) ? din_0_data[3] : wire_niiOliO_dataout;
	assign		wire_niiO0OO_dataout = (ni111ll === 1'b1) ? din_0_data[4] : wire_niiOlli_dataout;
	assign		wire_niiO10i_dataout = (ni111OO === 1'b1) ? niiiiOl : niii00i;
	assign		wire_niiO10l_dataout = (ni111OO === 1'b1) ? niiiiOO : niii00l;
	assign		wire_niiO10O_dataout = (ni111OO === 1'b1) ? niiil1i : niii00O;
	assign		wire_niiO11i_dataout = (ni111OO === 1'b1) ? niiiill : niii01i;
	assign		wire_niiO11l_dataout = (ni111OO === 1'b1) ? niiiilO : niii01l;
	assign		wire_niiO11O_dataout = (ni111OO === 1'b1) ? niiiiOi : niii01O;
	assign		wire_niiO1ii_dataout = (ni111OO === 1'b1) ? niiil1l : niii0ii;
	assign		wire_niiO1il_dataout = (ni111OO === 1'b1) ? niiil1O : niii0il;
	assign		wire_niiO1iO_dataout = (ni111OO === 1'b1) ? niiil0i : niii0iO;
	assign		wire_niiO1li_dataout = (ni111OO === 1'b1) ? niiil0l : niii0li;
	assign		wire_niiO1ll_dataout = (ni111OO === 1'b1) ? niiil0O : niii0ll;
	assign		wire_niiO1lO_dataout = (ni111OO === 1'b1) ? niiilii : niii0lO;
	assign		wire_niiO1Oi_dataout = (ni111OO === 1'b1) ? niiilil : niii0Oi;
	assign		wire_niiO1Ol_dataout = (ni111OO === 1'b1) ? niiiliO : niii0Ol;
	assign		wire_niiO1OO_dataout = (ni111OO === 1'b1) ? niiilli : niii0OO;
	assign		wire_niiOi0i_dataout = (ni111ll === 1'b1) ? din_0_data[8] : wire_niiOlOl_dataout;
	assign		wire_niiOi0l_dataout = (ni111ll === 1'b1) ? din_0_data[9] : wire_niiOlOO_dataout;
	assign		wire_niiOi0O_dataout = (ni111ll === 1'b1) ? din_0_data[10] : wire_niiOO1i_dataout;
	assign		wire_niiOi1i_dataout = (ni111ll === 1'b1) ? din_0_data[5] : wire_niiOlll_dataout;
	assign		wire_niiOi1l_dataout = (ni111ll === 1'b1) ? din_0_data[6] : wire_niiOllO_dataout;
	assign		wire_niiOi1O_dataout = (ni111ll === 1'b1) ? din_0_data[7] : wire_niiOlOi_dataout;
	assign		wire_niiOiii_dataout = (ni111ll === 1'b1) ? din_0_data[11] : wire_niiOO1l_dataout;
	assign		wire_niiOiil_dataout = (ni111ll === 1'b1) ? din_0_data[12] : wire_niiOO1O_dataout;
	assign		wire_niiOiiO_dataout = (ni111ll === 1'b1) ? din_0_data[13] : wire_niiOO0i_dataout;
	assign		wire_niiOili_dataout = (ni111ll === 1'b1) ? din_0_data[14] : wire_niiOO0l_dataout;
	assign		wire_niiOill_dataout = (ni111ll === 1'b1) ? din_0_data[15] : wire_niiOO0O_dataout;
	assign		wire_niiOilO_dataout = (ni111ll === 1'b1) ? din_0_data[16] : wire_niiOOii_dataout;
	assign		wire_niiOiOi_dataout = (ni111ll === 1'b1) ? din_0_data[17] : wire_niiOOil_dataout;
	assign		wire_niiOiOl_dataout = (ni111ll === 1'b1) ? din_0_data[18] : wire_niiOOiO_dataout;
	assign		wire_niiOiOO_dataout = (ni111ll === 1'b1) ? din_0_data[19] : wire_niiOOli_dataout;
	assign		wire_niiOl0i_dataout = (ni111ll === 1'b1) ? din_0_data[23] : wire_niiOOOl_dataout;
	assign		wire_niiOl0l_dataout = (ni111ll === 1'b1) ? din_0_endofpacket : wire_niiOOOO_dataout;
	assign		wire_niiOl0O_dataout = (ni111OO === 1'b1) ? niii1li : nii0lOO;
	assign		wire_niiOl1i_dataout = (ni111ll === 1'b1) ? din_0_data[20] : wire_niiOOll_dataout;
	assign		wire_niiOl1l_dataout = (ni111ll === 1'b1) ? din_0_data[21] : wire_niiOOlO_dataout;
	assign		wire_niiOl1O_dataout = (ni111ll === 1'b1) ? din_0_data[22] : wire_niiOOOi_dataout;
	assign		wire_niiOlii_dataout = (ni111OO === 1'b1) ? niii1ll : nii0O1i;
	assign		wire_niiOlil_dataout = (ni111OO === 1'b1) ? niii1lO : nii0O1l;
	assign		wire_niiOliO_dataout = (ni111OO === 1'b1) ? niii1Oi : nii0O1O;
	assign		wire_niiOlli_dataout = (ni111OO === 1'b1) ? niii1Ol : nii0O0i;
	assign		wire_niiOlll_dataout = (ni111OO === 1'b1) ? niii1OO : nii0O0l;
	assign		wire_niiOllO_dataout = (ni111OO === 1'b1) ? niii01i : nii0O0O;
	assign		wire_niiOlOi_dataout = (ni111OO === 1'b1) ? niii01l : nii0Oii;
	assign		wire_niiOlOl_dataout = (ni111OO === 1'b1) ? niii01O : nii0Oil;
	assign		wire_niiOlOO_dataout = (ni111OO === 1'b1) ? niii00i : nii0OiO;
	assign		wire_niiOO0i_dataout = (ni111OO === 1'b1) ? niii0il : nii0OOi;
	assign		wire_niiOO0l_dataout = (ni111OO === 1'b1) ? niii0iO : nii0OOl;
	assign		wire_niiOO0O_dataout = (ni111OO === 1'b1) ? niii0li : nii0OOO;
	assign		wire_niiOO1i_dataout = (ni111OO === 1'b1) ? niii00l : nii0Oli;
	assign		wire_niiOO1l_dataout = (ni111OO === 1'b1) ? niii00O : nii0Oll;
	assign		wire_niiOO1O_dataout = (ni111OO === 1'b1) ? niii0ii : nii0OlO;
	assign		wire_niiOOii_dataout = (ni111OO === 1'b1) ? niii0ll : niii11i;
	assign		wire_niiOOil_dataout = (ni111OO === 1'b1) ? niii0lO : niii11l;
	assign		wire_niiOOiO_dataout = (ni111OO === 1'b1) ? niii0Oi : niii11O;
	assign		wire_niiOOli_dataout = (ni111OO === 1'b1) ? niii0Ol : niii10i;
	assign		wire_niiOOll_dataout = (ni111OO === 1'b1) ? niii0OO : niii10l;
	assign		wire_niiOOlO_dataout = (ni111OO === 1'b1) ? niiii1i : niii10O;
	assign		wire_niiOOOi_dataout = (ni111OO === 1'b1) ? niiii1l : niii1ii;
	assign		wire_niiOOOl_dataout = (ni111OO === 1'b1) ? niiii1O : niii1il;
	assign		wire_niiOOOO_dataout = (ni111OO === 1'b1) ? niiii0i : niii1iO;
	and(wire_nil0O0i_dataout, nil1O1i, ~(ni110OO));
	assign		wire_nil0O0l_dataout = (ni110il === 1'b1) ? din_1_data[0] : wire_nili1OO_dataout;
	assign		wire_nil0O0O_dataout = (ni110il === 1'b1) ? din_1_data[1] : wire_nili01i_dataout;
	or(wire_nil0O1O_dataout, wire_nil0O0i_dataout, ni110il);
	assign		wire_nil0Oii_dataout = (ni110il === 1'b1) ? din_1_data[2] : wire_nili01l_dataout;
	assign		wire_nil0Oil_dataout = (ni110il === 1'b1) ? din_1_data[3] : wire_nili01O_dataout;
	assign		wire_nil0OiO_dataout = (ni110il === 1'b1) ? din_1_data[4] : wire_nili00i_dataout;
	assign		wire_nil0Oli_dataout = (ni110il === 1'b1) ? din_1_data[5] : wire_nili00l_dataout;
	assign		wire_nil0Oll_dataout = (ni110il === 1'b1) ? din_1_data[6] : wire_nili00O_dataout;
	assign		wire_nil0OlO_dataout = (ni110il === 1'b1) ? din_1_data[7] : wire_nili0ii_dataout;
	assign		wire_nil0OOi_dataout = (ni110il === 1'b1) ? din_1_data[8] : wire_nili0il_dataout;
	assign		wire_nil0OOl_dataout = (ni110il === 1'b1) ? din_1_data[9] : wire_nili0iO_dataout;
	assign		wire_nil0OOO_dataout = (ni110il === 1'b1) ? din_1_data[10] : wire_nili0li_dataout;
	and(wire_nil101i_dataout, nil11Ol, ~((~ ni1iili)));
	assign		wire_nil101l_dataout = ((~ ni1iili) === 1'b1) ? wire_nii00ii_o : nil11OO;
	assign		wire_nil10Oi_dataout = (nilO00l === 1'b1) ? wire_nil1i1i_dataout : wire_nil10Ol_dataout;
	or(wire_nil10Ol_dataout, wire_nil10OO_dataout, ni110Ol);
	assign		wire_nil10OO_dataout = (ni110Oi === 1'b1) ? (~ nil1lOO) : (~ nil1O1i);
	assign		wire_nil1i1i_dataout = (ni110Ol === 1'b1) ? (~ nil1O1i) : wire_nil1i1l_dataout;
	assign		wire_nil1i1l_dataout = (ni110Oi === 1'b1) ? (~ nil1lOi) : (~ nil1lOO);
	or(wire_nili00i_dataout, nil0ill, ni110OO);
	or(wire_nili00l_dataout, nil0ilO, ni110OO);
	or(wire_nili00O_dataout, nil0iOi, ni110OO);
	or(wire_nili01i_dataout, nil0iil, ni110OO);
	or(wire_nili01l_dataout, nil0iiO, ni110OO);
	or(wire_nili01O_dataout, nil0ili, ni110OO);
	or(wire_nili0ii_dataout, nil0iOl, ni110OO);
	or(wire_nili0il_dataout, nil0iOO, ni110OO);
	or(wire_nili0iO_dataout, nil0l1i, ni110OO);
	or(wire_nili0li_dataout, nil0l1l, ni110OO);
	or(wire_nili0ll_dataout, nil0l1O, ni110OO);
	or(wire_nili0lO_dataout, nil0l0i, ni110OO);
	or(wire_nili0Oi_dataout, nil0l0l, ni110OO);
	or(wire_nili0Ol_dataout, nil0l0O, ni110OO);
	or(wire_nili0OO_dataout, nil0lii, ni110OO);
	assign		wire_nili10i_dataout = (ni110il === 1'b1) ? din_1_data[14] : wire_nili0Ol_dataout;
	assign		wire_nili10l_dataout = (ni110il === 1'b1) ? din_1_data[15] : wire_nili0OO_dataout;
	assign		wire_nili10O_dataout = (ni110il === 1'b1) ? din_1_data[16] : wire_nilii1i_dataout;
	assign		wire_nili11i_dataout = (ni110il === 1'b1) ? din_1_data[11] : wire_nili0ll_dataout;
	assign		wire_nili11l_dataout = (ni110il === 1'b1) ? din_1_data[12] : wire_nili0lO_dataout;
	assign		wire_nili11O_dataout = (ni110il === 1'b1) ? din_1_data[13] : wire_nili0Oi_dataout;
	assign		wire_nili1ii_dataout = (ni110il === 1'b1) ? din_1_data[17] : wire_nilii1l_dataout;
	assign		wire_nili1il_dataout = (ni110il === 1'b1) ? din_1_data[18] : wire_nilii1O_dataout;
	assign		wire_nili1iO_dataout = (ni110il === 1'b1) ? din_1_data[19] : wire_nilii0i_dataout;
	assign		wire_nili1li_dataout = (ni110il === 1'b1) ? din_1_data[20] : wire_nilii0l_dataout;
	assign		wire_nili1ll_dataout = (ni110il === 1'b1) ? din_1_data[21] : wire_nilii0O_dataout;
	assign		wire_nili1lO_dataout = (ni110il === 1'b1) ? din_1_data[22] : wire_niliiii_dataout;
	assign		wire_nili1Oi_dataout = (ni110il === 1'b1) ? din_1_data[23] : wire_niliiil_dataout;
	assign		wire_nili1Ol_dataout = (ni110il === 1'b1) ? din_1_endofpacket : wire_niliiiO_dataout;
	or(wire_nili1OO_dataout, nil0iii, ni110OO);
	or(wire_nilii0i_dataout, nil0lll, ni110OO);
	or(wire_nilii0l_dataout, nil0llO, ni110OO);
	or(wire_nilii0O_dataout, nil0lOi, ni110OO);
	or(wire_nilii1i_dataout, nil0lil, ni110OO);
	or(wire_nilii1l_dataout, nil0liO, ni110OO);
	or(wire_nilii1O_dataout, nil0lli, ni110OO);
	or(wire_niliiii_dataout, nil0lOl, ni110OO);
	or(wire_niliiil_dataout, nil0lOO, ni110OO);
	or(wire_niliiiO_dataout, nil0O1i, ni110OO);
	or(wire_niliiOO_dataout, wire_nilil1i_dataout, ni110iO);
	assign		wire_nilil0i_dataout = (ni110iO === 1'b1) ? din_1_data[2] : wire_niliOOl_dataout;
	assign		wire_nilil0l_dataout = (ni110iO === 1'b1) ? din_1_data[3] : wire_niliOOO_dataout;
	assign		wire_nilil0O_dataout = (ni110iO === 1'b1) ? din_1_data[4] : wire_nill11i_dataout;
	assign		wire_nilil1i_dataout = (ni110OO === 1'b1) ? nil1O1i : nil1lOO;
	assign		wire_nilil1l_dataout = (ni110iO === 1'b1) ? din_1_data[0] : wire_niliOlO_dataout;
	assign		wire_nilil1O_dataout = (ni110iO === 1'b1) ? din_1_data[1] : wire_niliOOi_dataout;
	assign		wire_nililii_dataout = (ni110iO === 1'b1) ? din_1_data[5] : wire_nill11l_dataout;
	assign		wire_nililil_dataout = (ni110iO === 1'b1) ? din_1_data[6] : wire_nill11O_dataout;
	assign		wire_nililiO_dataout = (ni110iO === 1'b1) ? din_1_data[7] : wire_nill10i_dataout;
	assign		wire_nililli_dataout = (ni110iO === 1'b1) ? din_1_data[8] : wire_nill10l_dataout;
	assign		wire_nililll_dataout = (ni110iO === 1'b1) ? din_1_data[9] : wire_nill10O_dataout;
	assign		wire_nilillO_dataout = (ni110iO === 1'b1) ? din_1_data[10] : wire_nill1ii_dataout;
	assign		wire_nililOi_dataout = (ni110iO === 1'b1) ? din_1_data[11] : wire_nill1il_dataout;
	assign		wire_nililOl_dataout = (ni110iO === 1'b1) ? din_1_data[12] : wire_nill1iO_dataout;
	assign		wire_nililOO_dataout = (ni110iO === 1'b1) ? din_1_data[13] : wire_nill1li_dataout;
	assign		wire_niliO0i_dataout = (ni110iO === 1'b1) ? din_1_data[17] : wire_nill1Ol_dataout;
	assign		wire_niliO0l_dataout = (ni110iO === 1'b1) ? din_1_data[18] : wire_nill1OO_dataout;
	assign		wire_niliO0O_dataout = (ni110iO === 1'b1) ? din_1_data[19] : wire_nill01i_dataout;
	assign		wire_niliO1i_dataout = (ni110iO === 1'b1) ? din_1_data[14] : wire_nill1ll_dataout;
	assign		wire_niliO1l_dataout = (ni110iO === 1'b1) ? din_1_data[15] : wire_nill1lO_dataout;
	assign		wire_niliO1O_dataout = (ni110iO === 1'b1) ? din_1_data[16] : wire_nill1Oi_dataout;
	assign		wire_niliOii_dataout = (ni110iO === 1'b1) ? din_1_data[20] : wire_nill01l_dataout;
	assign		wire_niliOil_dataout = (ni110iO === 1'b1) ? din_1_data[21] : wire_nill01O_dataout;
	assign		wire_niliOiO_dataout = (ni110iO === 1'b1) ? din_1_data[22] : wire_nill00i_dataout;
	assign		wire_niliOli_dataout = (ni110iO === 1'b1) ? din_1_data[23] : wire_nill00l_dataout;
	assign		wire_niliOll_dataout = (ni110iO === 1'b1) ? din_1_endofpacket : wire_nill00O_dataout;
	assign		wire_niliOlO_dataout = (ni110OO === 1'b1) ? nil0iii : nil01lO;
	assign		wire_niliOOi_dataout = (ni110OO === 1'b1) ? nil0iil : nil01Oi;
	assign		wire_niliOOl_dataout = (ni110OO === 1'b1) ? nil0iiO : nil01Ol;
	assign		wire_niliOOO_dataout = (ni110OO === 1'b1) ? nil0ili : nil01OO;
	assign		wire_nill00i_dataout = (ni110OO === 1'b1) ? nil0lOl : nil0i0i;
	assign		wire_nill00l_dataout = (ni110OO === 1'b1) ? nil0lOO : nil0i0l;
	assign		wire_nill00O_dataout = (ni110OO === 1'b1) ? nil0O1i : nil0i0O;
	assign		wire_nill01i_dataout = (ni110OO === 1'b1) ? nil0lll : nil0i1i;
	assign		wire_nill01l_dataout = (ni110OO === 1'b1) ? nil0llO : nil0i1l;
	assign		wire_nill01O_dataout = (ni110OO === 1'b1) ? nil0lOi : nil0i1O;
	or(wire_nill0ll_dataout, wire_nill0lO_dataout, ni110ll);
	assign		wire_nill0lO_dataout = (ni110OO === 1'b1) ? nil1lOO : nil1lOi;
	assign		wire_nill0Oi_dataout = (ni110ll === 1'b1) ? din_1_data[0] : wire_nilllil_dataout;
	assign		wire_nill0Ol_dataout = (ni110ll === 1'b1) ? din_1_data[1] : wire_nillliO_dataout;
	assign		wire_nill0OO_dataout = (ni110ll === 1'b1) ? din_1_data[2] : wire_nilllli_dataout;
	assign		wire_nill10i_dataout = (ni110OO === 1'b1) ? nil0iOl : nil000i;
	assign		wire_nill10l_dataout = (ni110OO === 1'b1) ? nil0iOO : nil000l;
	assign		wire_nill10O_dataout = (ni110OO === 1'b1) ? nil0l1i : nil000O;
	assign		wire_nill11i_dataout = (ni110OO === 1'b1) ? nil0ill : nil001i;
	assign		wire_nill11l_dataout = (ni110OO === 1'b1) ? nil0ilO : nil001l;
	assign		wire_nill11O_dataout = (ni110OO === 1'b1) ? nil0iOi : nil001O;
	assign		wire_nill1ii_dataout = (ni110OO === 1'b1) ? nil0l1l : nil00ii;
	assign		wire_nill1il_dataout = (ni110OO === 1'b1) ? nil0l1O : nil00il;
	assign		wire_nill1iO_dataout = (ni110OO === 1'b1) ? nil0l0i : nil00iO;
	assign		wire_nill1li_dataout = (ni110OO === 1'b1) ? nil0l0l : nil00li;
	assign		wire_nill1ll_dataout = (ni110OO === 1'b1) ? nil0l0O : nil00ll;
	assign		wire_nill1lO_dataout = (ni110OO === 1'b1) ? nil0lii : nil00lO;
	assign		wire_nill1Oi_dataout = (ni110OO === 1'b1) ? nil0lil : nil00Oi;
	assign		wire_nill1Ol_dataout = (ni110OO === 1'b1) ? nil0liO : nil00Ol;
	assign		wire_nill1OO_dataout = (ni110OO === 1'b1) ? nil0lli : nil00OO;
	assign		wire_nilli0i_dataout = (ni110ll === 1'b1) ? din_1_data[6] : wire_nilllOl_dataout;
	assign		wire_nilli0l_dataout = (ni110ll === 1'b1) ? din_1_data[7] : wire_nilllOO_dataout;
	assign		wire_nilli0O_dataout = (ni110ll === 1'b1) ? din_1_data[8] : wire_nillO1i_dataout;
	assign		wire_nilli1i_dataout = (ni110ll === 1'b1) ? din_1_data[3] : wire_nilllll_dataout;
	assign		wire_nilli1l_dataout = (ni110ll === 1'b1) ? din_1_data[4] : wire_nillllO_dataout;
	assign		wire_nilli1O_dataout = (ni110ll === 1'b1) ? din_1_data[5] : wire_nilllOi_dataout;
	assign		wire_nilliii_dataout = (ni110ll === 1'b1) ? din_1_data[9] : wire_nillO1l_dataout;
	assign		wire_nilliil_dataout = (ni110ll === 1'b1) ? din_1_data[10] : wire_nillO1O_dataout;
	assign		wire_nilliiO_dataout = (ni110ll === 1'b1) ? din_1_data[11] : wire_nillO0i_dataout;
	assign		wire_nillili_dataout = (ni110ll === 1'b1) ? din_1_data[12] : wire_nillO0l_dataout;
	assign		wire_nillill_dataout = (ni110ll === 1'b1) ? din_1_data[13] : wire_nillO0O_dataout;
	assign		wire_nillilO_dataout = (ni110ll === 1'b1) ? din_1_data[14] : wire_nillOii_dataout;
	assign		wire_nilliOi_dataout = (ni110ll === 1'b1) ? din_1_data[15] : wire_nillOil_dataout;
	assign		wire_nilliOl_dataout = (ni110ll === 1'b1) ? din_1_data[16] : wire_nillOiO_dataout;
	assign		wire_nilliOO_dataout = (ni110ll === 1'b1) ? din_1_data[17] : wire_nillOli_dataout;
	assign		wire_nilll0i_dataout = (ni110ll === 1'b1) ? din_1_data[21] : wire_nillOOl_dataout;
	assign		wire_nilll0l_dataout = (ni110ll === 1'b1) ? din_1_data[22] : wire_nillOOO_dataout;
	assign		wire_nilll0O_dataout = (ni110ll === 1'b1) ? din_1_data[23] : wire_nilO11i_dataout;
	assign		wire_nilll1i_dataout = (ni110ll === 1'b1) ? din_1_data[18] : wire_nillOll_dataout;
	assign		wire_nilll1l_dataout = (ni110ll === 1'b1) ? din_1_data[19] : wire_nillOlO_dataout;
	assign		wire_nilll1O_dataout = (ni110ll === 1'b1) ? din_1_data[20] : wire_nillOOi_dataout;
	assign		wire_nilllii_dataout = (ni110ll === 1'b1) ? din_1_endofpacket : wire_nilO11l_dataout;
	assign		wire_nilllil_dataout = (ni110OO === 1'b1) ? nil01lO : nil1O1l;
	assign		wire_nillliO_dataout = (ni110OO === 1'b1) ? nil01Oi : nil1O1O;
	assign		wire_nilllli_dataout = (ni110OO === 1'b1) ? nil01Ol : nil1O0i;
	assign		wire_nilllll_dataout = (ni110OO === 1'b1) ? nil01OO : nil1O0l;
	assign		wire_nillllO_dataout = (ni110OO === 1'b1) ? nil001i : nil1O0O;
	assign		wire_nilllOi_dataout = (ni110OO === 1'b1) ? nil001l : nil1Oii;
	assign		wire_nilllOl_dataout = (ni110OO === 1'b1) ? nil001O : nil1Oil;
	assign		wire_nilllOO_dataout = (ni110OO === 1'b1) ? nil000i : nil1OiO;
	assign		wire_nillO0i_dataout = (ni110OO === 1'b1) ? nil00il : nil1OOi;
	assign		wire_nillO0l_dataout = (ni110OO === 1'b1) ? nil00iO : nil1OOl;
	assign		wire_nillO0O_dataout = (ni110OO === 1'b1) ? nil00li : nil1OOO;
	assign		wire_nillO1i_dataout = (ni110OO === 1'b1) ? nil000l : nil1Oli;
	assign		wire_nillO1l_dataout = (ni110OO === 1'b1) ? nil000O : nil1Oll;
	assign		wire_nillO1O_dataout = (ni110OO === 1'b1) ? nil00ii : nil1OlO;
	assign		wire_nillOii_dataout = (ni110OO === 1'b1) ? nil00ll : nil011i;
	assign		wire_nillOil_dataout = (ni110OO === 1'b1) ? nil00lO : nil011l;
	assign		wire_nillOiO_dataout = (ni110OO === 1'b1) ? nil00Oi : nil011O;
	assign		wire_nillOli_dataout = (ni110OO === 1'b1) ? nil00Ol : nil010i;
	assign		wire_nillOll_dataout = (ni110OO === 1'b1) ? nil00OO : nil010l;
	assign		wire_nillOlO_dataout = (ni110OO === 1'b1) ? nil0i1i : nil010O;
	assign		wire_nillOOi_dataout = (ni110OO === 1'b1) ? nil0i1l : nil01ii;
	assign		wire_nillOOl_dataout = (ni110OO === 1'b1) ? nil0i1O : nil01il;
	assign		wire_nillOOO_dataout = (ni110OO === 1'b1) ? nil0i0i : nil01iO;
	assign		wire_nilO00i_dataout = ((~ ni1iili) === 1'b1) ? wire_nil10iO_o : nilO01l;
	assign		wire_nilO00O_dataout = (nilOi0l === 1'b1) ? wire_nilO0il_dataout : wire_nilO0ii_dataout;
	and(wire_nilO01O_dataout, nilO01i, ~((~ ni1iili)));
	assign		wire_nilO0ii_dataout = (alpha_in_0_valid === 1'b1) ? (~ nilO0li) : (~ nilO0ll);
	assign		wire_nilO0il_dataout = (alpha_in_0_valid === 1'b1) ? (~ nilO0iO) : (~ nilO0li);
	or(wire_nilO0lO_dataout, nilO0ll, (alpha_in_0_valid & ((~ nilO0ll) & nilO0li)));
	or(wire_nilO0OO_dataout, nilO0li, (alpha_in_0_valid & ((~ nilO0li) & nilO0iO)));
	assign		wire_nilO11i_dataout = (ni110OO === 1'b1) ? nil0i0l : nil01li;
	assign		wire_nilO11l_dataout = (ni110OO === 1'b1) ? nil0i0O : nil01ll;
	or(wire_nilOi1l_dataout, nilO0iO, (alpha_in_0_valid & (~ nilO0iO)));
	assign		wire_nilOiOO_dataout = (niO00lO === 1'b1) ? wire_nilOl1O_dataout : wire_nilOl1i_dataout;
	assign		wire_nilOl0i_dataout = (ni11iOi === 1'b1) ? (~ nilOlOl) : (~ nilOO1i);
	or(wire_nilOl1i_dataout, wire_nilOl1l_dataout, ni11iOl);
	assign		wire_nilOl1l_dataout = (ni11iOi === 1'b1) ? (~ nilOO1i) : (~ nilOO1l);
	assign		wire_nilOl1O_dataout = (ni11iOl === 1'b1) ? (~ nilOO1l) : wire_nilOl0i_dataout;
	and(wire_niO00li_dataout, niO00il, ~((~ ni1iili)));
	assign		wire_niO00ll_dataout = ((~ ni1iili) === 1'b1) ? wire_nilOill_o : niO00iO;
	assign		wire_niO010i_dataout = (ni11iOO === 1'b1) ? nilOOOO : nilOO0O;
	assign		wire_niO010l_dataout = (ni11iOO === 1'b1) ? niO111i : nilOOii;
	assign		wire_niO010O_dataout = (ni11iOO === 1'b1) ? niO111l : nilOOil;
	assign		wire_niO011i_dataout = (ni11iOO === 1'b1) ? nilOOlO : nilOO1O;
	assign		wire_niO011l_dataout = (ni11iOO === 1'b1) ? nilOOOi : nilOO0i;
	assign		wire_niO011O_dataout = (ni11iOO === 1'b1) ? nilOOOl : nilOO0l;
	assign		wire_niO01ii_dataout = (ni11iOO === 1'b1) ? niO111O : nilOOiO;
	assign		wire_niO01il_dataout = (ni11iOO === 1'b1) ? niO110i : nilOOli;
	assign		wire_niO01iO_dataout = (ni11iOO === 1'b1) ? niO110l : nilOOll;
	assign		wire_niO100i_dataout = (ni11iil === 1'b1) ? alpha_in_1_data[1] : wire_niO10Oi_dataout;
	assign		wire_niO100l_dataout = (ni11iil === 1'b1) ? alpha_in_1_data[2] : wire_niO10Ol_dataout;
	assign		wire_niO100O_dataout = (ni11iil === 1'b1) ? alpha_in_1_data[3] : wire_niO10OO_dataout;
	or(wire_niO101i_dataout, wire_niO101l_dataout, ni11iil);
	and(wire_niO101l_dataout, nilOO1l, ~(ni11iOO));
	assign		wire_niO101O_dataout = (ni11iil === 1'b1) ? alpha_in_1_data[0] : wire_niO10lO_dataout;
	assign		wire_niO10ii_dataout = (ni11iil === 1'b1) ? alpha_in_1_data[4] : wire_niO1i1i_dataout;
	assign		wire_niO10il_dataout = (ni11iil === 1'b1) ? alpha_in_1_data[5] : wire_niO1i1l_dataout;
	assign		wire_niO10iO_dataout = (ni11iil === 1'b1) ? alpha_in_1_data[6] : wire_niO1i1O_dataout;
	assign		wire_niO10li_dataout = (ni11iil === 1'b1) ? alpha_in_1_data[7] : wire_niO1i0i_dataout;
	assign		wire_niO10ll_dataout = (ni11iil === 1'b1) ? alpha_in_1_endofpacket : wire_niO1i0l_dataout;
	or(wire_niO10lO_dataout, niO110O, ni11iOO);
	or(wire_niO10Oi_dataout, niO11ii, ni11iOO);
	or(wire_niO10Ol_dataout, niO11il, ni11iOO);
	or(wire_niO10OO_dataout, niO11iO, ni11iOO);
	or(wire_niO1i0i_dataout, niO11Oi, ni11iOO);
	or(wire_niO1i0l_dataout, niO11Ol, ni11iOO);
	or(wire_niO1i1i_dataout, niO11li, ni11iOO);
	or(wire_niO1i1l_dataout, niO11ll, ni11iOO);
	or(wire_niO1i1O_dataout, niO11lO, ni11iOO);
	or(wire_niO1ill_dataout, wire_niO1ilO_dataout, ni11iiO);
	assign		wire_niO1ilO_dataout = (ni11iOO === 1'b1) ? nilOO1l : nilOO1i;
	assign		wire_niO1iOi_dataout = (ni11iiO === 1'b1) ? alpha_in_1_data[0] : wire_niO1lii_dataout;
	assign		wire_niO1iOl_dataout = (ni11iiO === 1'b1) ? alpha_in_1_data[1] : wire_niO1lil_dataout;
	assign		wire_niO1iOO_dataout = (ni11iiO === 1'b1) ? alpha_in_1_data[2] : wire_niO1liO_dataout;
	assign		wire_niO1l0i_dataout = (ni11iiO === 1'b1) ? alpha_in_1_data[6] : wire_niO1lOi_dataout;
	assign		wire_niO1l0l_dataout = (ni11iiO === 1'b1) ? alpha_in_1_data[7] : wire_niO1lOl_dataout;
	assign		wire_niO1l0O_dataout = (ni11iiO === 1'b1) ? alpha_in_1_endofpacket : wire_niO1lOO_dataout;
	assign		wire_niO1l1i_dataout = (ni11iiO === 1'b1) ? alpha_in_1_data[3] : wire_niO1lli_dataout;
	assign		wire_niO1l1l_dataout = (ni11iiO === 1'b1) ? alpha_in_1_data[4] : wire_niO1lll_dataout;
	assign		wire_niO1l1O_dataout = (ni11iiO === 1'b1) ? alpha_in_1_data[5] : wire_niO1llO_dataout;
	assign		wire_niO1lii_dataout = (ni11iOO === 1'b1) ? niO110O : nilOOlO;
	assign		wire_niO1lil_dataout = (ni11iOO === 1'b1) ? niO11ii : nilOOOi;
	assign		wire_niO1liO_dataout = (ni11iOO === 1'b1) ? niO11il : nilOOOl;
	assign		wire_niO1lli_dataout = (ni11iOO === 1'b1) ? niO11iO : nilOOOO;
	assign		wire_niO1lll_dataout = (ni11iOO === 1'b1) ? niO11li : niO111i;
	assign		wire_niO1llO_dataout = (ni11iOO === 1'b1) ? niO11ll : niO111l;
	assign		wire_niO1lOi_dataout = (ni11iOO === 1'b1) ? niO11lO : niO111O;
	assign		wire_niO1lOl_dataout = (ni11iOO === 1'b1) ? niO11Oi : niO110i;
	assign		wire_niO1lOO_dataout = (ni11iOO === 1'b1) ? niO11Ol : niO110l;
	or(wire_niO1O0l_dataout, wire_niO1O0O_dataout, ni11ill);
	assign		wire_niO1O0O_dataout = (ni11iOO === 1'b1) ? nilOO1i : nilOlOl;
	assign		wire_niO1Oii_dataout = (ni11ill === 1'b1) ? alpha_in_1_data[0] : wire_niO011i_dataout;
	assign		wire_niO1Oil_dataout = (ni11ill === 1'b1) ? alpha_in_1_data[1] : wire_niO011l_dataout;
	assign		wire_niO1OiO_dataout = (ni11ill === 1'b1) ? alpha_in_1_data[2] : wire_niO011O_dataout;
	assign		wire_niO1Oli_dataout = (ni11ill === 1'b1) ? alpha_in_1_data[3] : wire_niO010i_dataout;
	assign		wire_niO1Oll_dataout = (ni11ill === 1'b1) ? alpha_in_1_data[4] : wire_niO010l_dataout;
	assign		wire_niO1OlO_dataout = (ni11ill === 1'b1) ? alpha_in_1_data[5] : wire_niO010O_dataout;
	assign		wire_niO1OOi_dataout = (ni11ill === 1'b1) ? alpha_in_1_data[6] : wire_niO01ii_dataout;
	assign		wire_niO1OOl_dataout = (ni11ill === 1'b1) ? alpha_in_1_data[7] : wire_niO01il_dataout;
	assign		wire_niO1OOO_dataout = (ni11ill === 1'b1) ? alpha_in_1_endofpacket : wire_niO01iO_dataout;
	and(wire_niOiOil_dataout, wire_niOiOiO_dataout, ~(dout_ready));
	or(wire_niOiOiO_dataout, niOii0l, ((~ dout_ready) & ni11Oii));
	and(wire_niOl00i_dataout, nl00OOl, ~(ni11Oli));
	and(wire_niOl00l_dataout, nl00OOO, ~(ni11Oli));
	and(wire_niOl00O_dataout, nl0i11i, ~(ni11Oli));
	assign		wire_niOl01i_dataout = (ni11OiO === 1'b1) ? nl00lil : wire_niOl0ii_dataout;
	and(wire_niOl01l_dataout, nl00OlO, ~(ni11Oli));
	and(wire_niOl01O_dataout, nl00OOi, ~(ni11Oli));
	and(wire_niOl0ii_dataout, nl0i11O, ~(ni11Oli));
	assign		wire_niOl10l_dataout = (ni11Oil === 1'b1) ? n0Oll : wire_niOl1ll_dataout;
	and(wire_niOl10O_dataout, wire_niOl1lO_dataout, ~(ni11Oil));
	and(wire_niOl1ii_dataout, wire_niOl1Oi_dataout, ~(ni11Oil));
	and(wire_niOl1il_dataout, wire_niOl1Ol_dataout, ~(ni11Oil));
	and(wire_niOl1iO_dataout, wire_niOl1OO_dataout, ~(ni11Oil));
	and(wire_niOl1li_dataout, wire_niOl01i_dataout, ~(ni11Oil));
	assign		wire_niOl1ll_dataout = (ni11OiO === 1'b1) ? nl00l1l : wire_niOl01l_dataout;
	assign		wire_niOl1lO_dataout = (ni11OiO === 1'b1) ? nl00l1O : wire_niOl01O_dataout;
	assign		wire_niOl1Oi_dataout = (ni11OiO === 1'b1) ? nl00l0i : wire_niOl00i_dataout;
	assign		wire_niOl1Ol_dataout = (ni11OiO === 1'b1) ? nl00l0l : wire_niOl00l_dataout;
	assign		wire_niOl1OO_dataout = (ni11OiO === 1'b1) ? nl00l0O : wire_niOl00O_dataout;
	and(wire_nl0i00i_dataout, wire_nl0i0il_o[5], ~(n0Oll));
	and(wire_nl0i00l_dataout, wire_nl0i0il_o[6], ~(n0Oll));
	and(wire_nl0i00O_dataout, wire_nl0i0il_o[7], ~(n0Oll));
	and(wire_nl0i01i_dataout, wire_nl0i0il_o[2], ~(n0Oll));
	and(wire_nl0i01l_dataout, wire_nl0i0il_o[3], ~(n0Oll));
	and(wire_nl0i01O_dataout, wire_nl0i0il_o[4], ~(n0Oll));
	and(wire_nl0i0ii_dataout, wire_nl0i0il_o[8], ~(n0Oll));
	and(wire_nl0i1OO_dataout, wire_nl0i0il_o[1], ~(n0Oll));
	and(wire_nl0iill_dataout, wire_nl0il0O_o[1], ~(n00ii));
	and(wire_nl0iilO_dataout, wire_nl0il0O_o[2], ~(n00ii));
	and(wire_nl0iiOi_dataout, wire_nl0il0O_o[3], ~(n00ii));
	and(wire_nl0iiOl_dataout, wire_nl0il0O_o[4], ~(n00ii));
	and(wire_nl0iiOO_dataout, wire_nl0il0O_o[5], ~(n00ii));
	and(wire_nl0il0i_dataout, wire_nl0il0O_o[9], ~(n00ii));
	and(wire_nl0il0l_dataout, wire_nl0il0O_o[10], ~(n00ii));
	and(wire_nl0il1i_dataout, wire_nl0il0O_o[6], ~(n00ii));
	and(wire_nl0il1l_dataout, wire_nl0il0O_o[7], ~(n00ii));
	and(wire_nl0il1O_dataout, wire_nl0il0O_o[8], ~(n00ii));
	and(wire_nl0iO0i_dataout, wire_nl0iOOl_o[1], ~(n00ii));
	and(wire_nl0iO0l_dataout, wire_nl0iOOl_o[2], ~(n00ii));
	and(wire_nl0iO0O_dataout, wire_nl0iOOl_o[3], ~(n00ii));
	and(wire_nl0iOii_dataout, wire_nl0iOOl_o[4], ~(n00ii));
	and(wire_nl0iOil_dataout, wire_nl0iOOl_o[5], ~(n00ii));
	and(wire_nl0iOiO_dataout, wire_nl0iOOl_o[6], ~(n00ii));
	and(wire_nl0iOli_dataout, wire_nl0iOOl_o[7], ~(n00ii));
	and(wire_nl0iOll_dataout, wire_nl0iOOl_o[8], ~(n00ii));
	and(wire_nl0iOlO_dataout, wire_nl0iOOl_o[9], ~(n00ii));
	and(wire_nl0iOOi_dataout, wire_nl0iOOl_o[10], ~(n00ii));
	or(wire_nl0l01i_dataout, wire_nl0l01O_o[2], n11ll);
	and(wire_nl0l01l_dataout, wire_nl0l01O_o[3], ~(n11ll));
	assign		wire_nl0O10i_dataout = ((~ n11li) === 1'b1) ? wire_nl0O1Oi_o[4] : wire_nl0O1lO_o[5];
	assign		wire_nl0O10l_dataout = ((~ n11li) === 1'b1) ? wire_nl0O1Oi_o[5] : wire_nl0O1lO_o[6];
	assign		wire_nl0O10O_dataout = ((~ n11li) === 1'b1) ? wire_nl0O1Oi_o[6] : wire_nl0O1lO_o[7];
	assign		wire_nl0O11i_dataout = ((~ n11li) === 1'b1) ? wire_nl0O1Oi_o[1] : wire_nl0O1lO_o[2];
	assign		wire_nl0O11l_dataout = ((~ n11li) === 1'b1) ? wire_nl0O1Oi_o[2] : wire_nl0O1lO_o[3];
	assign		wire_nl0O11O_dataout = ((~ n11li) === 1'b1) ? wire_nl0O1Oi_o[3] : wire_nl0O1lO_o[4];
	assign		wire_nl0O1ii_dataout = ((~ n11li) === 1'b1) ? wire_nl0O1Oi_o[7] : wire_nl0O1lO_o[8];
	assign		wire_nl0O1il_dataout = ((~ n11li) === 1'b1) ? wire_nl0O1Oi_o[8] : wire_nl0O1lO_o[9];
	assign		wire_nl0O1iO_dataout = ((~ n11li) === 1'b1) ? wire_nl0O1Oi_o[9] : wire_nl0O1lO_o[10];
	assign		wire_nl0O1li_dataout = ((~ n11li) === 1'b1) ? wire_nl0O1Oi_o[10] : wire_nl0O1lO_o[11];
	assign		wire_nl0O1ll_dataout = ((~ n11li) === 1'b1) ? wire_nl0O1Oi_o[11] : wire_nl0O1lO_o[12];
	assign		wire_nl1lO0l_dataout = (wire_nl1lliO_o === 1'b1) ? wire_nl1liOi_o : wire_nl1lOOi_o[1];
	assign		wire_nl1lO0O_dataout = (wire_nl1lliO_o === 1'b1) ? wire_nl1liOl_o : wire_nl1lOOi_o[2];
	assign		wire_nl1lOii_dataout = (wire_nl1lliO_o === 1'b1) ? wire_nl1liOO_o : wire_nl1lOOi_o[3];
	assign		wire_nl1lOil_dataout = (wire_nl1lliO_o === 1'b1) ? wire_nl1ll1i_o : wire_nl1lOOi_o[4];
	assign		wire_nl1lOiO_dataout = (wire_nl1lliO_o === 1'b1) ? wire_nl1ll1l_o : wire_nl1lOOi_o[5];
	assign		wire_nl1lOli_dataout = (wire_nl1lliO_o === 1'b1) ? wire_nl1ll1O_o : wire_nl1lOOi_o[6];
	assign		wire_nl1lOll_dataout = (wire_nl1lliO_o === 1'b1) ? wire_nl1ll0i_o : wire_nl1lOOi_o[7];
	assign		wire_nl1lOlO_dataout = (wire_nl1lliO_o === 1'b1) ? wire_nl1ll0l_o : wire_nl1lOOi_o[8];
	and(wire_nl1O0ii_dataout, wire_nl1Oi1i_o[2], ~(ni1i10i));
	and(wire_nl1O0il_dataout, wire_nl1Oi1i_o[3], ~(ni1i10i));
	and(wire_nl1O0iO_dataout, wire_nl1Oi1i_o[4], ~(ni1i10i));
	and(wire_nl1O0li_dataout, wire_nl1Oi1i_o[5], ~(ni1i10i));
	and(wire_nl1O0ll_dataout, wire_nl1Oi1i_o[6], ~(ni1i10i));
	and(wire_nl1O0lO_dataout, wire_nl1Oi1i_o[7], ~(ni1i10i));
	and(wire_nl1O0Oi_dataout, wire_nl1Oi1i_o[8], ~(ni1i10i));
	and(wire_nl1O0Ol_dataout, wire_nl1Oi1i_o[9], ~(ni1i10i));
	and(wire_nl1O0OO_dataout, wire_nl1Oi1i_o[10], ~(ni1i10i));
	oper_add   ni010Ol
	( 
	.a({ni0100l, ni01i1O}),
	.b({1'b0, 1'b1}),
	.cin(1'b0),
	.cout(),
	.o(wire_ni010Ol_o));
	defparam
		ni010Ol.sgate_representation = 0,
		ni010Ol.width_a = 2,
		ni010Ol.width_b = 2,
		ni010Ol.width_o = 2;
	oper_add   ni01i1l
	( 
	.a({ni0100l, ni01i1O, 1'b1}),
	.b({1'b1, 1'b0, 1'b1}),
	.cin(1'b0),
	.cout(),
	.o(wire_ni01i1l_o));
	defparam
		ni01i1l.sgate_representation = 0,
		ni01i1l.width_a = 3,
		ni01i1l.width_b = 3,
		ni01i1l.width_o = 3;
	oper_add   ni01iOO
	( 
	.a({ni01iii, ni010ii}),
	.b({1'b0, 1'b1}),
	.cin(1'b0),
	.cout(),
	.o(wire_ni01iOO_o));
	defparam
		ni01iOO.sgate_representation = 0,
		ni01iOO.width_a = 2,
		ni01iOO.width_b = 2,
		ni01iOO.width_o = 2;
	oper_add   ni01l0i
	( 
	.a({ni01iii, ni010ii, 1'b1}),
	.b({1'b1, 1'b0, 1'b1}),
	.cin(1'b0),
	.cout(),
	.o(wire_ni01l0i_o));
	defparam
		ni01l0i.sgate_representation = 0,
		ni01l0i.width_a = 3,
		ni01l0i.width_b = 3,
		ni01l0i.width_o = 3;
	oper_add   ni01lOO
	( 
	.a({ni01lli, ni01liO}),
	.b({1'b0, 1'b1}),
	.cin(1'b0),
	.cout(),
	.o(wire_ni01lOO_o));
	defparam
		ni01lOO.sgate_representation = 0,
		ni01lOO.width_a = 2,
		ni01lOO.width_b = 2,
		ni01lOO.width_o = 2;
	oper_add   ni01O1O
	( 
	.a({ni01lli, ni01liO, 1'b1}),
	.b({1'b1, 1'b0, 1'b1}),
	.cin(1'b0),
	.cout(),
	.o(wire_ni01O1O_o));
	defparam
		ni01O1O.sgate_representation = 0,
		ni01O1O.width_a = 3,
		ni01O1O.width_b = 3,
		ni01O1O.width_o = 3;
	oper_add   ni0Oiil
	( 
	.a({ni0Oi1O}),
	.b({1'b1}),
	.cin(1'b0),
	.cout(),
	.o(wire_ni0Oiil_o));
	defparam
		ni0Oiil.sgate_representation = 0,
		ni0Oiil.width_a = 1,
		ni0Oiil.width_b = 1,
		ni0Oiil.width_o = 1;
	oper_add   ni0Oili
	( 
	.a({ni0Oi1O, 1'b1}),
	.b({1'b0, 1'b1}),
	.cin(1'b0),
	.cout(),
	.o(wire_ni0Oili_o));
	defparam
		ni0Oili.sgate_representation = 0,
		ni0Oili.width_a = 2,
		ni0Oili.width_b = 2,
		ni0Oili.width_o = 2;
	oper_add   nii001l
	( 
	.a({nii01il, nii01ii, nii010O, nii010l, nii010i, nii01li, 1'b0}),
	.b({{4{1'b0}}, n0Oil, 1'b1, 1'b0}),
	.cin(1'b0),
	.cout(),
	.o(wire_nii001l_o));
	defparam
		nii001l.sgate_representation = 0,
		nii001l.width_a = 7,
		nii001l.width_b = 7,
		nii001l.width_o = 7;
	oper_add   nii011l
	( 
	.a({nii1Oli, nii1OiO, nii1Oil, nii1OlO, 1'b0}),
	.b({{3{1'b0}}, 1'b1, 1'b0}),
	.cin(1'b0),
	.cout(),
	.o(wire_nii011l_o));
	defparam
		nii011l.sgate_representation = 0,
		nii011l.width_a = 5,
		nii011l.width_b = 5,
		nii011l.width_o = 5;
	oper_add   niOO1lO
	( 
	.a({niOliil, niOliii, niOli0O, niOli0l, niOli0i, niOli1O, niOli1l, niOli1i, niOl0OO, niOlili, 1'b0}),
	.b({nl1i11i, nl10OOl, nl10OlO, nl10Oll, nl10Oli, nl10OiO, nl10Oil, nl10Oii, nl10O0O, nl10O0l, 1'b0}),
	.cin(1'b0),
	.cout(),
	.o(wire_niOO1lO_o));
	defparam
		niOO1lO.sgate_representation = 0,
		niOO1lO.width_a = 11,
		niOO1lO.width_b = 11,
		niOO1lO.width_o = 11;
	oper_add   niOOi0l
	( 
	.a({niOO0ii, niOO00l, niOO00i, niOO01O, niOO01l, niOO01i, niOO1OO, niOO1Ol, 1'b0}),
	.b({nl1i0li, nl1i0il, nl1i0ii, nl1i00O, nl1i00l, nl1i01O, nl1i01l, nl1i01i, 1'b0}),
	.cin(1'b0),
	.cout(),
	.o(wire_niOOi0l_o));
	defparam
		niOOi0l.sgate_representation = 0,
		niOOi0l.width_a = 9,
		niOOi0l.width_b = 9,
		niOOi0l.width_o = 9;
	oper_add   nl0i0il
	( 
	.a({nl0i1lO, nl0i1ll, nl0i1li, nl0i1iO, nl0i1il, nl0i1ii, nl0i10O, nl0i1Ol, 1'b0}),
	.b({{7{1'b0}}, 1'b1, 1'b0}),
	.cin(1'b0),
	.cout(),
	.o(wire_nl0i0il_o));
	defparam
		nl0i0il.sgate_representation = 0,
		nl0i0il.width_a = 9,
		nl0i0il.width_b = 9,
		nl0i0il.width_o = 9;
	oper_add   nl0il0O
	( 
	.a({nl0iiil, nl0iiii, nl0ii0O, nl0ii0l, nl0ii0i, nl0ii1O, nl0ii1l, nl0ii1i, nl0i0OO, nl0iili, 1'b0}),
	.b({{9{1'b0}}, 1'b1, 1'b0}),
	.cin(1'b0),
	.cout(),
	.o(wire_nl0il0O_o));
	defparam
		nl0il0O.sgate_representation = 0,
		nl0il0O.width_a = 11,
		nl0il0O.width_b = 11,
		nl0il0O.width_o = 11;
	oper_add   nl0iOOl
	( 
	.a({nl0iO1i, nl0ilOO, nl0ilOl, nl0ilOi, nl0illO, nl0illl, nl0illi, nl0iliO, nl0ilil, nl0iO1O, 1'b0}),
	.b({{9{1'b0}}, 1'b1, 1'b0}),
	.cin(1'b0),
	.cout(),
	.o(wire_nl0iOOl_o));
	defparam
		nl0iOOl.sgate_representation = 0,
		nl0iOOl.width_a = 11,
		nl0iOOl.width_b = 11,
		nl0iOOl.width_o = 11;
	oper_add   nl0l01O
	( 
	.a({nl0l1Oi, nl0l1OO, 1'b0, 1'b1}),
	.b({1'b1, 1'b0, {2{1'b1}}}),
	.cin(1'b0),
	.cout(),
	.o(wire_nl0l01O_o));
	defparam
		nl0l01O.sgate_representation = 0,
		nl0l01O.width_a = 4,
		nl0l01O.width_b = 4,
		nl0l01O.width_o = 4;
	oper_add   nl0O00O
	( 
	.a({1'b0, nl0i1lO, nl0i1ll, nl0i1li, nl0i1iO, nl0i1il, nl0i1ii, nl0i10O, nl0i1Ol, 1'b1}),
	.b({1'b1, (~ nl1i1Oi), (~ nl1i1ll), (~ nl1i1li), (~ nl1i1iO), (~ nl1i1il), (~ nl1i10O), (~ nl1i10l), (~ nl1i10i), 1'b1}),
	.cin(1'b0),
	.cout(),
	.o(wire_nl0O00O_o));
	defparam
		nl0O00O.sgate_representation = 0,
		nl0O00O.width_a = 10,
		nl0O00O.width_b = 10,
		nl0O00O.width_o = 10;
	oper_add   nl0O0ii
	( 
	.a({1'b0, nl0iO1i, nl0ilOO, nl0ilOl, nl0ilOi, nl0illO, nl0illl, nl0illi, nl0iliO, nl0ilil, nl0iO1O, 1'b1}),
	.b({1'b1, (~ niOlOli), (~ niOlOiO), (~ niOlOil), (~ niOlOii), (~ niOlO0O), (~ niOlO0l), (~ niOlO0i), (~ niOlO1O), (~ niOlO1l), (~ niOlOlO), 1'b1}),
	.cin(1'b0),
	.cout(),
	.o(wire_nl0O0ii_o));
	defparam
		nl0O0ii.sgate_representation = 0,
		nl0O0ii.width_a = 12,
		nl0O0ii.width_b = 12,
		nl0O0ii.width_o = 12;
	oper_add   nl0O1lO
	( 
	.a({wire_nl0lO1l_o, wire_nl0lO1i_o, wire_nl0llOO_o, wire_nl0llOl_o, wire_nl0llOi_o, wire_nl0lllO_o, wire_nl0llll_o, wire_nl0llli_o, wire_nl0lliO_o, wire_nl0llil_o, wire_nl0llii_o, 1'b0, 1'b1}),
	.b({{10{(~ n111l)}}, 1'b0, {2{1'b1}}}),
	.cin(1'b0),
	.cout(),
	.o(wire_nl0O1lO_o));
	defparam
		nl0O1lO.sgate_representation = 0,
		nl0O1lO.width_a = 13,
		nl0O1lO.width_b = 13,
		nl0O1lO.width_o = 13;
	oper_add   nl0O1Oi
	( 
	.a({wire_nl0lO1l_o, wire_nl0lO1i_o, wire_nl0llOO_o, wire_nl0llOl_o, wire_nl0llOi_o, wire_nl0lllO_o, wire_nl0llll_o, wire_nl0llli_o, wire_nl0lliO_o, wire_nl0llil_o, wire_nl0llii_o, 1'b0}),
	.b({{10{n111l}}, 1'b1, 1'b0}),
	.cin(1'b0),
	.cout(),
	.o(wire_nl0O1Oi_o));
	defparam
		nl0O1Oi.sgate_representation = 0,
		nl0O1Oi.width_a = 12,
		nl0O1Oi.width_b = 12,
		nl0O1Oi.width_o = 12;
	oper_add   nl0Olil
	( 
	.a({nl1i1Oi, nl1i1ll, nl1i1li, nl1i1iO, nl1i1il, nl1i10O, nl1i10l, nl1i10i, 1'b0}),
	.b({{8{1'b1}}, 1'b0}),
	.cin(1'b0),
	.cout(),
	.o(wire_nl0Olil_o));
	defparam
		nl0Olil.sgate_representation = 0,
		nl0Olil.width_a = 9,
		nl0Olil.width_b = 9,
		nl0Olil.width_o = 9;
	oper_add   nl0OOii
	( 
	.a({1'b0, nl0iiil, nl0iiii, nl0ii0O, nl0ii0l, nl0ii0i, nl0ii1O, nl0ii1l, nl0ii1i, nl0i0OO, nl0iili, 1'b1}),
	.b({1'b1, (~ niOliil), (~ niOliii), (~ niOli0O), (~ niOli0l), (~ niOli0i), (~ niOli1O), (~ niOli1l), (~ niOli1i), (~ niOl0OO), (~ niOlili), 1'b1}),
	.cin(1'b0),
	.cout(),
	.o(wire_nl0OOii_o));
	defparam
		nl0OOii.sgate_representation = 0,
		nl0OOii.width_a = 12,
		nl0OOii.width_b = 12,
		nl0OOii.width_o = 12;
	oper_add   nl1iOll
	( 
	.a({1'b0, wire_nl1Oi1O_result[16:0], 1'b0}),
	.b({1'b0, wire_nl1Ol0O_result[16:0], 1'b0}),
	.cin(1'b0),
	.cout(),
	.o(wire_nl1iOll_o));
	defparam
		nl1iOll.sgate_representation = 0,
		nl1iOll.width_a = 19,
		nl1iOll.width_b = 19,
		nl1iOll.width_o = 19;
	oper_add   nl1l01O
	( 
	.a({1'b0, wire_nl1OiOO_result[16:0], 1'b0}),
	.b({1'b0, wire_nl1OO1O_result[16:0], 1'b0}),
	.cin(1'b0),
	.cout(),
	.o(wire_nl1l01O_o));
	defparam
		nl1l01O.sgate_representation = 0,
		nl1l01O.width_a = 19,
		nl1l01O.width_b = 19,
		nl1l01O.width_o = 19;
	oper_add   nl1l1ii
	( 
	.a({1'b0, wire_nl1OiiO_result[16:0], 1'b0}),
	.b({1'b0, wire_nl1OllO_result[16:0], 1'b0}),
	.cin(1'b0),
	.cout(),
	.o(wire_nl1l1ii_o));
	defparam
		nl1l1ii.sgate_representation = 0,
		nl1l1ii.width_a = 19,
		nl1l1ii.width_b = 19,
		nl1l1ii.width_o = 19;
	oper_add   nl1lOOi
	( 
	.a({wire_nl1li0i_o, wire_nl1li1O_o, wire_nl1li1l_o, wire_nl1li1i_o, wire_nl1l0OO_o, wire_nl1l0Ol_o, wire_nl1l0Oi_o, wire_nl1l0lO_o, 1'b0}),
	.b({9{1'b0}}),
	.cin(1'b0),
	.cout(),
	.o(wire_nl1lOOi_o));
	defparam
		nl1lOOi.sgate_representation = 0,
		nl1lOOi.width_a = 9,
		nl1lOOi.width_b = 9,
		nl1lOOi.width_o = 9;
	oper_add   nl1Oi1i
	( 
	.a({1'b1, (~ nl1lO1l), (~ nl1lO1i), (~ nl1llOO), (~ nl1llOl), (~ nl1llOi), (~ nl1lllO), (~ nl1llll), (~ nl1lO0i), {2{1'b1}}}),
	.b({1'b1, {9{1'b0}}, 1'b1}),
	.cin(1'b0),
	.cout(),
	.o(wire_nl1Oi1i_o));
	defparam
		nl1Oi1i.sgate_representation = 0,
		nl1Oi1i.width_a = 11,
		nl1Oi1i.width_b = 11,
		nl1Oi1i.width_o = 11;
	oper_add   nli110l
	( 
	.a({1'b0, nl0iiil, nl0iiii, nl0ii0O, nl0ii0l, nl0ii0i, nl0ii1O, nl0ii1l, nl0ii1i, nl0i0OO, nl0iili, 1'b1}),
	.b({1'b1, (~ niOO1iO), (~ niOO1il), (~ niOO1ii), (~ niOO10O), (~ niOO10l), (~ niOO10i), (~ niOO11O), (~ niOO11l), (~ niOO11i), (~ niOO1ll), 1'b1}),
	.cin(1'b0),
	.cout(),
	.o(wire_nli110l_o));
	defparam
		nli110l.sgate_representation = 0,
		nli110l.width_a = 12,
		nli110l.width_b = 12,
		nli110l.width_o = 12;
	oper_add   nli110O
	( 
	.a({1'b0, nl0i1lO, nl0i1ll, nl0i1li, nl0i1iO, nl0i1il, nl0i1ii, nl0i10O, nl0i1Ol, 1'b1}),
	.b({1'b1, (~ niOO0ii), (~ niOO00l), (~ niOO00i), (~ niOO01O), (~ niOO01l), (~ niOO01i), (~ niOO1OO), (~ niOO1Ol), 1'b1}),
	.cin(1'b0),
	.cout(),
	.o(wire_nli110O_o));
	defparam
		nli110O.sgate_representation = 0,
		nli110O.width_a = 10,
		nli110O.width_b = 10,
		nli110O.width_o = 10;
	oper_add   nli11ii
	( 
	.a({1'b0, nl0i1lO, nl0i1ll, nl0i1li, nl0i1iO, nl0i1il, nl0i1ii, nl0i10O, nl0i1Ol, 1'b1}),
	.b({1'b1, (~ niOOi1l), (~ niOOi1i), (~ niOO0OO), (~ niOO0Ol), (~ niOO0Oi), (~ niOO0lO), (~ niOO0ll), (~ niOOi0i), 1'b1}),
	.cin(1'b0),
	.cout(),
	.o(wire_nli11ii_o));
	defparam
		nli11ii.sgate_representation = 0,
		nli11ii.width_a = 10,
		nli11ii.width_b = 10,
		nli11ii.width_o = 10;
	oper_less_than   nii111l
	( 
	.a({1'b0}),
	.b({ni0Oi1O}),
	.cin(1'b0),
	.o(wire_nii111l_o));
	defparam
		nii111l.sgate_representation = 0,
		nii111l.width_a = 1,
		nii111l.width_b = 1;
	oper_mux   n011i
	( 
	.data({{76{ni1iOli}}, 1'b1, {42{1'b0}}, 1'b1, {8{1'b0}}}),
	.o(wire_n011i_o),
	.sel({n1ili, n1iil, n1iii, n1i0O, n1i0l, n1i0i, n1i1O}));
	defparam
		n011i.width_data = 128,
		n011i.width_sel = 7;
	oper_mux   n011l
	( 
	.data({{108{ni1iOli}}, 1'b1, {11{1'b0}}, 1'b1, {7{1'b0}}}),
	.o(wire_n011l_o),
	.sel({n1ili, n1iil, n1iii, n1i0O, n1i0l, n1i0i, n1i1O}));
	defparam
		n011l.width_data = 128,
		n011l.width_sel = 7;
	oper_mux   n1ilO
	( 
	.data({{3{1'b0}}, 1'b1}),
	.o(wire_n1ilO_o),
	.sel({n1i0l, n1i0i}));
	defparam
		n1ilO.width_data = 4,
		n1ilO.width_sel = 2;
	oper_mux   n1iOi
	( 
	.data({{9{1'b0}}, 1'b1, {5{1'b0}}, 1'b1}),
	.o(wire_n1iOi_o),
	.sel({n1ili, n1i0l, n1i0i, n1i1O}));
	defparam
		n1iOi.width_data = 16,
		n1iOi.width_sel = 4;
	oper_mux   n1iOl
	( 
	.data({{3{1'b0}}, 1'b1, {4{1'b0}}, 1'b1, {4{1'b0}}, 1'b1, {2{1'b0}}}),
	.o(wire_n1iOl_o),
	.sel({n1i0O, n1i0l, n1i0i, n1i1O}));
	defparam
		n1iOl.width_data = 16,
		n1iOl.width_sel = 4;
	oper_mux   n1iOO
	( 
	.data({{13{1'b0}}, 1'b1, {10{1'b0}}, {6{1'b1}}, {3{1'b0}}, 1'b1, {30{1'b0}}}),
	.o(wire_n1iOO_o),
	.sel({n1iil, n1iii, n1i0O, n1i0l, n1i0i, n1i1O}));
	defparam
		n1iOO.width_data = 64,
		n1iOO.width_sel = 6;
	oper_mux   n1l0i
	( 
	.data({1'b0, 1'b1, {6{1'b0}}, 1'b1, {2{1'b0}}, 1'b1, 1'b0, 1'b1, {2{1'b0}}}),
	.o(wire_n1l0i_o),
	.sel({n1iil, n1i0O, n1i0l, n1i0i}));
	defparam
		n1l0i.width_data = 16,
		n1l0i.width_sel = 4;
	oper_mux   n1l0l
	( 
	.data({{3{1'b0}}, 1'b1, {5{1'b0}}, 1'b1, {5{1'b0}}, 1'b1}),
	.o(wire_n1l0l_o),
	.sel({n1ili, n1i0O, n1i0l, n1i0i}));
	defparam
		n1l0l.width_data = 16,
		n1l0l.width_sel = 4;
	oper_mux   n1l0O
	( 
	.data({{2{1'b0}}, {2{1'b1}}, {3{1'b0}}, {2{1'b1}}, {3{1'b0}}, 1'b1, {8{1'b0}}, {5{1'b1}}, {6{1'b0}}, 1'b1, {17{1'b0}}, {2{1'b1}}, {2{1'b0}}, 1'b1, {3{1'b0}}, 1'b1, {3{1'b0}}, 1'b1, 1'b0}),
	.o(wire_n1l0O_o),
	.sel({n1iil, n1iii, n1i0O, n1i0l, n1i0i, n1i1O}));
	defparam
		n1l0O.width_data = 64,
		n1l0O.width_sel = 6;
	oper_mux   n1l1i
	( 
	.data({{5{1'b1}}, {2{1'b0}}, 1'b1}),
	.o(wire_n1l1i_o),
	.sel({n1iii, n1i0O, n1i0l}));
	defparam
		n1l1i.width_data = 8,
		n1l1i.width_sel = 3;
	oper_mux   n1l1l
	( 
	.data({{3{1'b0}}, 1'b1, {5{1'b0}}, 1'b1, {3{1'b0}}, 1'b1, 1'b0, 1'b1}),
	.o(wire_n1l1l_o),
	.sel({n1iil, n1iii, n1i0O, n1i1O}));
	defparam
		n1l1l.width_data = 16,
		n1l1l.width_sel = 4;
	oper_mux   n1l1O
	( 
	.data({{11{ni1iOli}}, 1'b1, {9{1'b0}}, {5{1'b1}}, {6{1'b0}}}),
	.o(wire_n1l1O_o),
	.sel({n1ili, n1i0O, n1i0l, n1i0i, n1i1O}));
	defparam
		n1l1O.width_data = 32,
		n1l1O.width_sel = 5;
	oper_mux   n1lii
	( 
	.data({{15{ni1iOli}}, 1'b1}),
	.o(wire_n1lii_o),
	.sel({n1ili, n1iii, n1i0i, n1i1O}));
	defparam
		n1lii.width_data = 16,
		n1lii.width_sel = 4;
	oper_mux   n1lil
	( 
	.data({{86{ni1iOli}}, {5{1'b1}}, {11{1'b0}}, 1'b1, {13{1'b0}}, 1'b1, {4{1'b0}}, 1'b1, {6{1'b0}}}),
	.o(wire_n1lil_o),
	.sel({n1ili, n1iil, n1iii, n1i0O, n1i0l, n1i0i, n1i1O}));
	defparam
		n1lil.width_data = 128,
		n1lil.width_sel = 7;
	oper_mux   n1liO
	( 
	.data({{4{1'b0}}, 1'b1, {4{1'b0}}, 1'b1, {53{1'b0}}, 1'b1}),
	.o(wire_n1liO_o),
	.sel({n1iil, n1iii, n1i0O, n1i0l, n1i0i, n1i1O}));
	defparam
		n1liO.width_data = 64,
		n1liO.width_sel = 6;
	oper_mux   n1lli
	( 
	.data({{84{ni1iOli}}, {10{1'b1}}, {14{1'b0}}, 1'b1, {15{1'b0}}, 1'b1, {3{1'b0}}}),
	.o(wire_n1lli_o),
	.sel({n1ili, n1iil, n1iii, n1i0O, n1i0l, n1i0i, n1i1O}));
	defparam
		n1lli.width_data = 128,
		n1lli.width_sel = 7;
	oper_mux   n1lll
	( 
	.data({{55{ni1iOli}}, 1'b1, {63{1'b0}}, 1'b1, {4{1'b0}}, 1'b1, {3{1'b0}}}),
	.o(wire_n1lll_o),
	.sel({n1ili, n1iil, n1iii, n1i0O, n1i0l, n1i0i, n1i1O}));
	defparam
		n1lll.width_data = 128,
		n1lll.width_sel = 7;
	oper_mux   n1llO
	( 
	.data({{54{ni1iOli}}, 1'b1, {45{1'b0}}, 1'b1, {27{1'b0}}}),
	.o(wire_n1llO_o),
	.sel({n1ili, n1iil, n1iii, n1i0O, n1i0l, n1i0i, n1i1O}));
	defparam
		n1llO.width_data = 128,
		n1llO.width_sel = 7;
	oper_mux   n1lOi
	( 
	.data({{53{ni1iOli}}, 1'b1, {30{1'b0}}, {5{1'b1}}, {11{1'b0}}, 1'b1, {27{1'b0}}}),
	.o(wire_n1lOi_o),
	.sel({n1ili, n1iil, n1iii, n1i0O, n1i0l, n1i0i, n1i1O}));
	defparam
		n1lOi.width_data = 128,
		n1lOi.width_sel = 7;
	oper_mux   n1lOl
	( 
	.data({{12{1'b0}}, 1'b1, {51{1'b0}}}),
	.o(wire_n1lOl_o),
	.sel({n1iil, n1iii, n1i0O, n1i0l, n1i0i, n1i1O}));
	defparam
		n1lOl.width_data = 64,
		n1lOl.width_sel = 6;
	oper_mux   n1lOO
	( 
	.data({{62{ni1iOli}}, 1'b1, {4{1'b0}}, 1'b1, {4{1'b0}}, 1'b1, {55{1'b0}}}),
	.o(wire_n1lOO_o),
	.sel({n1ili, n1iil, n1iii, n1i0O, n1i0l, n1i0i, n1i1O}));
	defparam
		n1lOO.width_data = 128,
		n1lOO.width_sel = 7;
	oper_mux   n1O0i
	( 
	.data({{19{1'b0}}, 1'b1, {44{1'b0}}}),
	.o(wire_n1O0i_o),
	.sel({n1iil, n1iii, n1i0O, n1i0l, n1i0i, n1i1O}));
	defparam
		n1O0i.width_data = 64,
		n1O0i.width_sel = 6;
	oper_mux   n1O0l
	( 
	.data({{43{1'b0}}, 1'b1, {20{1'b0}}}),
	.o(wire_n1O0l_o),
	.sel({n1iil, n1iii, n1i0O, n1i0l, n1i0i, n1i1O}));
	defparam
		n1O0l.width_data = 64,
		n1O0l.width_sel = 6;
	oper_mux   n1O0O
	( 
	.data({{14{ni1iOli}}, 1'b1, {17{1'b0}}}),
	.o(wire_n1O0O_o),
	.sel({n1ili, n1i0O, n1i0l, n1i0i, n1i1O}));
	defparam
		n1O0O.width_data = 32,
		n1O0O.width_sel = 5;
	oper_mux   n1O1i
	( 
	.data({{51{ni1iOli}}, 1'b1, {28{1'b0}}, 1'b1, {47{1'b0}}}),
	.o(wire_n1O1i_o),
	.sel({n1ili, n1iil, n1iii, n1i0O, n1i0l, n1i0i, n1i1O}));
	defparam
		n1O1i.width_data = 128,
		n1O1i.width_sel = 7;
	oper_mux   n1O1l
	( 
	.data({{36{1'b0}}, 1'b1, {27{1'b0}}}),
	.o(wire_n1O1l_o),
	.sel({n1iil, n1iii, n1i0O, n1i0l, n1i0i, n1i1O}));
	defparam
		n1O1l.width_data = 64,
		n1O1l.width_sel = 6;
	oper_mux   n1O1O
	( 
	.data({{32{1'b0}}, 1'b1, {31{1'b0}}}),
	.o(wire_n1O1O_o),
	.sel({n1iil, n1iii, n1i0O, n1i0l, n1i0i, n1i1O}));
	defparam
		n1O1O.width_data = 64,
		n1O1O.width_sel = 6;
	oper_mux   n1Oii
	( 
	.data({{6{ni1iOli}}, 1'b1, {25{1'b0}}}),
	.o(wire_n1Oii_o),
	.sel({n1ili, n1i0O, n1i0l, n1i0i, n1i1O}));
	defparam
		n1Oii.width_data = 32,
		n1Oii.width_sel = 5;
	oper_mux   n1Oil
	( 
	.data({{111{ni1iOli}}, 1'b1, {2{1'b0}}, 1'b1, {13{1'b0}}}),
	.o(wire_n1Oil_o),
	.sel({n1ili, n1iil, n1iii, n1i0O, n1i0l, n1i0i, n1i1O}));
	defparam
		n1Oil.width_data = 128,
		n1Oil.width_sel = 7;
	oper_mux   n1OiO
	( 
	.data({{88{ni1iOli}}, {5{1'b1}}, {11{1'b0}}, 1'b1, {13{1'b0}}, 1'b1, {4{1'b0}}, 1'b1, {4{1'b0}}}),
	.o(wire_n1OiO_o),
	.sel({n1ili, n1iil, n1iii, n1i0O, n1i0l, n1i0i, n1i1O}));
	defparam
		n1OiO.width_data = 128,
		n1OiO.width_sel = 7;
	oper_mux   n1Oli
	( 
	.data({1'b0, 1'b1, {4{1'b0}}, 1'b1, {4{1'b0}}, 1'b1, {52{1'b0}}}),
	.o(wire_n1Oli_o),
	.sel({n1iil, n1iii, n1i0O, n1i0l, n1i0i, n1i1O}));
	defparam
		n1Oli.width_data = 64,
		n1Oli.width_sel = 6;
	oper_mux   n1Oll
	( 
	.data({{9{ni1iOli}}, 1'b1, {22{1'b0}}}),
	.o(wire_n1Oll_o),
	.sel({n1ili, n1i0O, n1i0l, n1i0i, n1i1O}));
	defparam
		n1Oll.width_data = 32,
		n1Oll.width_sel = 5;
	oper_mux   n1OlO
	( 
	.data({{12{ni1iOli}}, 1'b1, {19{1'b0}}}),
	.o(wire_n1OlO_o),
	.sel({n1ili, n1i0O, n1i0l, n1i0i, n1i1O}));
	defparam
		n1OlO.width_data = 32,
		n1OlO.width_sel = 5;
	oper_mux   n1OOi
	( 
	.data({{2{1'b0}}, 1'b1, {61{1'b0}}}),
	.o(wire_n1OOi_o),
	.sel({n1iil, n1iii, n1i0O, n1i0l, n1i0i, n1i1O}));
	defparam
		n1OOi.width_data = 64,
		n1OOi.width_sel = 6;
	oper_mux   n1OOl
	( 
	.data({{24{1'b0}}, 1'b1, {39{1'b0}}}),
	.o(wire_n1OOl_o),
	.sel({n1iil, n1iii, n1i0O, n1i0l, n1i0i, n1i1O}));
	defparam
		n1OOl.width_data = 64,
		n1OOl.width_sel = 6;
	oper_mux   n1OOO
	( 
	.data({{53{ni1iOli}}, 1'b1, {8{1'b0}}, 1'b1, {4{1'b0}}, 1'b1, {4{1'b0}}, 1'b1, {3{1'b0}}, 1'b1, {6{1'b0}}, {6{1'b1}}, {11{1'b0}}, 1'b1, {27{1'b0}}}),
	.o(wire_n1OOO_o),
	.sel({n1ili, n1iil, n1iii, n1i0O, n1i0l, n1i0i, n1i1O}));
	defparam
		n1OOO.width_data = 128,
		n1OOO.width_sel = 7;
	oper_mux   ni00i
	( 
	.data({{30{ni1iOli}}, 1'b1, {3{1'b0}}, {2{1'b1}}, {8{1'b0}}, 1'b1, {4{1'b0}}, 1'b1, {2{1'b0}}, {5{1'b1}}, {2{1'b0}}, 1'b1, {3{1'b0}}, 1'b1}),
	.o(wire_ni00i_o),
	.sel({ni10l, ni11O, ni11l, ni11i, n0OOO, n0OOi}));
	defparam
		ni00i.width_data = 64,
		ni00i.width_sel = 6;
	oper_mux   ni00l
	( 
	.data({{31{ni1iOli}}, 1'b1, 1'b0, {2{1'b1}}, {10{1'b0}}, 1'b1, {2{1'b0}}, 1'b1, {2{1'b0}}, 1'b1, 1'b0, 1'b1, 1'b0, {2{1'b1}}, {3{1'b0}}, 1'b1, {3{1'b0}}}),
	.o(wire_ni00l_o),
	.sel({ni10l, ni11O, ni11l, n0OOO, n0OOl, n0OOi}));
	defparam
		ni00l.width_data = 64,
		ni00l.width_sel = 6;
	oper_mux   ni00O
	( 
	.data({{30{ni1iOli}}, 1'b1, {6{1'b0}}, {2{1'b1}}, {2{1'b0}}, 1'b1, {8{1'b0}}, 1'b1, 1'b0, 1'b1, {2{1'b0}}, {2{1'b1}}, 1'b0, 1'b1, {5{1'b0}}}),
	.o(wire_ni00O_o),
	.sel({ni10l, ni11l, ni11i, n0OOO, n0OOl, n0OOi}));
	defparam
		ni00O.width_data = 64,
		ni00O.width_sel = 6;
	oper_mux   ni01i
	( 
	.data({{7{1'b0}}, {2{1'b1}}, {7{1'b0}}}),
	.o(wire_ni01i_o),
	.sel({n0OOO, n0OOl, n0OOi, n0OlO}));
	defparam
		ni01i.width_data = 16,
		ni01i.width_sel = 4;
	oper_mux   ni01l
	( 
	.data({{47{1'b0}}, 1'b1, {12{1'b0}}, 1'b1, {3{1'b0}}}),
	.o(wire_ni01l_o),
	.sel({ni11O, ni11l, ni11i, n0OOO, n0OOl, n0OOi}));
	defparam
		ni01l.width_data = 64,
		ni01l.width_sel = 6;
	oper_mux   ni01O
	( 
	.data({1'b1, 1'b0, {2{1'b1}}, {13{1'b0}}, 1'b1, 1'b0, 1'b1, 1'b0, {2{1'b1}}, {3{1'b0}}, {2{1'b1}}, {3{1'b0}}, 1'b1}),
	.o(wire_ni01O_o),
	.sel({ni11O, ni11l, ni11i, n0OOO, n0OOi}));
	defparam
		ni01O.width_data = 32,
		ni01O.width_sel = 5;
	oper_mux   ni0ii
	( 
	.data({{15{ni1iOli}}, {3{1'b1}}, {2{1'b0}}, {2{1'b1}}, 1'b0, 1'b1, {8{1'b0}}}),
	.o(wire_ni0ii_o),
	.sel({ni10l, ni11O, ni11l, n0OOO, n0OOi}));
	defparam
		ni0ii.width_data = 32,
		ni0ii.width_sel = 5;
	oper_mux   ni0il
	( 
	.data({{43{ni1iOli}}, 1'b1, {9{1'b0}}, {2{1'b1}}, {4{1'b0}}, {2{1'b1}}, {3{1'b0}}}),
	.o(wire_ni0il_o),
	.sel({ni10l, ni11O, ni11l, ni11i, n0OOi, n0OlO}));
	defparam
		ni0il.width_data = 64,
		ni0il.width_sel = 6;
	oper_mux   ni0iO
	( 
	.data({1'b0, 1'b1, {2{1'b0}}}),
	.o(wire_ni0iO_o),
	.sel({ni11i, n0OOl}));
	defparam
		ni0iO.width_data = 4,
		ni0iO.width_sel = 2;
	oper_mux   ni0li
	( 
	.data({{16{ni1iOli}}, {2{1'b1}}, {3{1'b0}}, {3{1'b1}}, {2{1'b0}}, 1'b1, {2{1'b0}}, 1'b1, 1'b0, 1'b1}),
	.o(wire_ni0li_o),
	.sel({ni10l, ni11O, ni11i, n0OOO, n0OOl}));
	defparam
		ni0li.width_data = 32,
		ni0li.width_sel = 5;
	oper_mux   ni0ll
	( 
	.data({{124{ni1iOli}}, 1'b1, {45{1'b0}}, {2{1'b1}}, {2{1'b0}}, 1'b1, {6{1'b0}}, 1'b1, {20{1'b0}}, 1'b1, {2{1'b0}}, 1'b1, {2{1'b0}}, {3{1'b1}}, {3{1'b0}}, 1'b1, {5{1'b0}}, 1'b1, {2{1'b0}}, 1'b1, {2{1'b0}}, 1'b1, {15{1'b0}}, {2{1'b1}}, {12{1'b0}}}),
	.o(wire_ni0ll_o),
	.sel({ni10l, ni11O, ni11l, ni11i, n0OOO, n0OOl, n0OOi, n0OlO}));
	defparam
		ni0ll.width_data = 256,
		ni0ll.width_sel = 8;
	oper_mux   ni0lO
	( 
	.data({{147{ni1iOli}}, 1'b1, {27{1'b0}}, 1'b1, {6{1'b0}}, 1'b1, {8{1'b0}}, 1'b1, {60{1'b0}}, 1'b1, {3{1'b0}}}),
	.o(wire_ni0lO_o),
	.sel({ni10l, ni11O, ni11l, ni11i, n0OOO, n0OOl, n0OOi, n0OlO}));
	defparam
		ni0lO.width_data = 256,
		ni0lO.width_sel = 8;
	oper_mux   ni0Oi
	( 
	.data({1'b0, {2{1'b1}}, {125{1'b0}}}),
	.o(wire_ni0Oi_o),
	.sel({ni11O, ni11l, ni11i, n0OOO, n0OOl, n0OOi, n0OlO}));
	defparam
		ni0Oi.width_data = 128,
		ni0Oi.width_sel = 7;
	oper_mux   ni0Ol
	( 
	.data({{55{1'b0}}, 1'b1, {72{1'b0}}}),
	.o(wire_ni0Ol_o),
	.sel({ni11O, ni11l, ni11i, n0OOO, n0OOl, n0OOi, n0OlO}));
	defparam
		ni0Ol.width_data = 128,
		ni0Ol.width_sel = 7;
	oper_mux   ni0OO
	( 
	.data({{27{1'b0}}, {10{1'b1}}, {91{1'b0}}}),
	.o(wire_ni0OO_o),
	.sel({ni11O, ni11l, ni11i, n0OOO, n0OOl, n0OOi, n0OlO}));
	defparam
		ni0OO.width_data = 128,
		ni0OO.width_sel = 7;
	oper_mux   ni10O
	( 
	.data({{9{ni1iOli}}, {7{1'b1}}}),
	.o(wire_ni10O_o),
	.sel({ni10l, n0OOO, n0OOi, n0OlO}));
	defparam
		ni10O.width_data = 16,
		ni10O.width_sel = 4;
	oper_mux   ni1ii
	( 
	.data({{5{ni1iOli}}, {3{1'b1}}}),
	.o(wire_ni1ii_o),
	.sel({ni10l, n0OOO, n0OOi}));
	defparam
		ni1ii.width_data = 8,
		ni1ii.width_sel = 3;
	oper_mux   ni1il
	( 
	.data({1'b0, {4{1'b1}}, {3{1'b0}}}),
	.o(wire_ni1il_o),
	.sel({ni11l, n0OOO, n0OlO}));
	defparam
		ni1il.width_data = 8,
		ni1il.width_sel = 3;
	oper_mux   ni1iO
	( 
	.data({1'b0, {2{1'b1}}, 1'b0}),
	.o(wire_ni1iO_o),
	.sel({ni11l, n0OOO}));
	defparam
		ni1iO.width_data = 4,
		ni1iO.width_sel = 2;
	oper_mux   ni1li
	( 
	.data({{17{ni1iOli}}, {10{1'b1}}, {5{1'b0}}}),
	.o(wire_ni1li_o),
	.sel({ni10l, ni11l, n0OOl, n0OOi, n0OlO}));
	defparam
		ni1li.width_data = 32,
		ni1li.width_sel = 5;
	oper_mux   ni1ll
	( 
	.data({{45{ni1iOli}}, {11{1'b1}}, {3{1'b0}}, 1'b1, {4{1'b0}}}),
	.o(wire_ni1ll_o),
	.sel({ni10l, ni11l, n0OOO, n0OOl, n0OOi, n0OlO}));
	defparam
		ni1ll.width_data = 64,
		ni1ll.width_sel = 6;
	oper_mux   ni1lO
	( 
	.data({{45{ni1iOli}}, {10{1'b1}}, {4{1'b0}}, 1'b1, {4{1'b0}}}),
	.o(wire_ni1lO_o),
	.sel({ni10l, ni11l, n0OOO, n0OOl, n0OOi, n0OlO}));
	defparam
		ni1lO.width_data = 64,
		ni1lO.width_sel = 6;
	oper_mux   ni1Oi
	( 
	.data({{13{1'b0}}, {5{1'b1}}, {9{1'b0}}, 1'b1, {4{1'b0}}}),
	.o(wire_ni1Oi_o),
	.sel({ni11l, ni11i, n0OOO, n0OOl, n0OOi}));
	defparam
		ni1Oi.width_data = 32,
		ni1Oi.width_sel = 5;
	oper_mux   ni1Ol
	( 
	.data({{3{1'b0}}, 1'b1}),
	.o(wire_ni1Ol_o),
	.sel({ni10l, n0OOl}));
	defparam
		ni1Ol.width_data = 4,
		ni1Ol.width_sel = 2;
	oper_mux   ni1OO
	( 
	.data({{8{ni1iOli}}, {4{1'b1}}, {3{1'b0}}, 1'b1}),
	.o(wire_ni1OO_o),
	.sel({ni10l, ni11O, n0OOO, n0OlO}));
	defparam
		ni1OO.width_data = 16,
		ni1OO.width_sel = 4;
	oper_mux   nii0i
	( 
	.data({{29{1'b0}}, 1'b1, {98{1'b0}}}),
	.o(wire_nii0i_o),
	.sel({ni11O, ni11l, ni11i, n0OOO, n0OOl, n0OOi, n0OlO}));
	defparam
		nii0i.width_data = 128,
		nii0i.width_sel = 7;
	oper_mux   nii0l
	( 
	.data({{109{1'b0}}, 1'b1, {18{1'b0}}}),
	.o(wire_nii0l_o),
	.sel({ni11O, ni11l, ni11i, n0OOO, n0OOl, n0OOi, n0OlO}));
	defparam
		nii0l.width_data = 128,
		nii0l.width_sel = 7;
	oper_mux   nii0O
	( 
	.data({1'b0, 1'b1, {126{1'b0}}}),
	.o(wire_nii0O_o),
	.sel({ni11O, ni11l, ni11i, n0OOO, n0OOl, n0OOi, n0OlO}));
	defparam
		nii0O.width_data = 128,
		nii0O.width_sel = 7;
	oper_mux   nii1i
	( 
	.data({{5{1'b0}}, 1'b1, {58{1'b0}}}),
	.o(wire_nii1i_o),
	.sel({ni11O, ni11l, ni11i, n0OOO, n0OOl, n0OOi}));
	defparam
		nii1i.width_data = 64,
		nii1i.width_sel = 6;
	oper_mux   nii1l
	( 
	.data({{41{1'b0}}, 1'b1, {22{1'b0}}}),
	.o(wire_nii1l_o),
	.sel({ni11O, ni11l, ni11i, n0OOO, n0OOl, n0OOi}));
	defparam
		nii1l.width_data = 64,
		nii1l.width_sel = 6;
	oper_mux   nii1O
	( 
	.data({{89{1'b0}}, 1'b1, {38{1'b0}}}),
	.o(wire_nii1O_o),
	.sel({ni11O, ni11l, ni11i, n0OOO, n0OOl, n0OOi, n0OlO}));
	defparam
		nii1O.width_data = 128,
		nii1O.width_sel = 7;
	oper_mux   niiii
	( 
	.data({{10{1'b0}}, 1'b1, {117{1'b0}}}),
	.o(wire_niiii_o),
	.sel({ni11O, ni11l, ni11i, n0OOO, n0OOl, n0OOi, n0OlO}));
	defparam
		niiii.width_data = 128,
		niiii.width_sel = 7;
	oper_mux   niiil
	( 
	.data({{82{1'b0}}, 1'b1, {45{1'b0}}}),
	.o(wire_niiil_o),
	.sel({ni11O, ni11l, ni11i, n0OOO, n0OOl, n0OOi, n0OlO}));
	defparam
		niiil.width_data = 128,
		niiil.width_sel = 7;
	oper_mux   niiiO
	( 
	.data({{10{1'b0}}, {2{1'b1}}, {17{1'b0}}, {10{1'b1}}, {70{1'b0}}, {2{1'b1}}, {17{1'b0}}}),
	.o(wire_niiiO_o),
	.sel({ni11O, ni11l, ni11i, n0OOO, n0OOl, n0OOi, n0OlO}));
	defparam
		niiiO.width_data = 128,
		niiiO.width_sel = 7;
	oper_mux   niili
	( 
	.data({{116{1'b0}}, 1'b1, {11{1'b0}}}),
	.o(wire_niili_o),
	.sel({ni11O, ni11l, ni11i, n0OOO, n0OOl, n0OOi, n0OlO}));
	defparam
		niili.width_data = 128,
		niili.width_sel = 7;
	oper_mux   niill
	( 
	.data({{124{ni1iOli}}, 1'b1, {2{1'b0}}, 1'b1, {8{1'b0}}, 1'b1, {119{1'b0}}}),
	.o(wire_niill_o),
	.sel({ni10l, ni11O, ni11l, ni11i, n0OOO, n0OOl, n0OOi, n0OlO}));
	defparam
		niill.width_data = 256,
		niill.width_sel = 8;
	oper_mux   niilO
	( 
	.data({{14{1'b0}}, 1'b1, {113{1'b0}}}),
	.o(wire_niilO_o),
	.sel({ni11O, ni11l, ni11i, n0OOO, n0OOl, n0OOi, n0OlO}));
	defparam
		niilO.width_data = 128,
		niilO.width_sel = 7;
	oper_mux   niiOi
	( 
	.data({{107{1'b0}}, 1'b1, {20{1'b0}}}),
	.o(wire_niiOi_o),
	.sel({ni11O, ni11l, ni11i, n0OOO, n0OOl, n0OOi, n0OlO}));
	defparam
		niiOi.width_data = 128,
		niiOi.width_sel = 7;
	oper_mux   niiOl
	( 
	.data({{80{1'b0}}, 1'b1, {47{1'b0}}}),
	.o(wire_niiOl_o),
	.sel({ni11O, ni11l, ni11i, n0OOO, n0OOl, n0OOi, n0OlO}));
	defparam
		niiOl.width_data = 128,
		niiOl.width_sel = 7;
	oper_mux   niiOO
	( 
	.data({{66{1'b0}}, 1'b1, {61{1'b0}}}),
	.o(wire_niiOO_o),
	.sel({ni11O, ni11l, ni11i, n0OOO, n0OOl, n0OOi, n0OlO}));
	defparam
		niiOO.width_data = 128,
		niiOO.width_sel = 7;
	oper_mux   nil0i
	( 
	.data({{46{1'b0}}, 1'b1, {81{1'b0}}}),
	.o(wire_nil0i_o),
	.sel({ni11O, ni11l, ni11i, n0OOO, n0OOl, n0OOi, n0OlO}));
	defparam
		nil0i.width_data = 128,
		nil0i.width_sel = 7;
	oper_mux   nil0l
	( 
	.data({{42{1'b0}}, 1'b1, {85{1'b0}}}),
	.o(wire_nil0l_o),
	.sel({ni11O, ni11l, ni11i, n0OOO, n0OOl, n0OOi, n0OlO}));
	defparam
		nil0l.width_data = 128,
		nil0l.width_sel = 7;
	oper_mux   nil0O
	( 
	.data({{18{1'b0}}, 1'b1, {109{1'b0}}}),
	.o(wire_nil0O_o),
	.sel({ni11O, ni11l, ni11i, n0OOO, n0OOl, n0OOi, n0OlO}));
	defparam
		nil0O.width_data = 128,
		nil0O.width_sel = 7;
	oper_mux   nil1i
	( 
	.data({{50{1'b0}}, 1'b1, {2{1'b0}}, 1'b1, {74{1'b0}}}),
	.o(wire_nil1i_o),
	.sel({ni11O, ni11l, ni11i, n0OOO, n0OOl, n0OOi, n0OlO}));
	defparam
		nil1i.width_data = 128,
		nil1i.width_sel = 7;
	oper_mux   nil1l
	( 
	.data({{113{1'b0}}, 1'b1, {14{1'b0}}}),
	.o(wire_nil1l_o),
	.sel({ni11O, ni11l, ni11i, n0OOO, n0OOl, n0OOi, n0OlO}));
	defparam
		nil1l.width_data = 128,
		nil1l.width_sel = 7;
	oper_mux   nil1O
	( 
	.data({{5{1'b0}}, 1'b1, {122{1'b0}}}),
	.o(wire_nil1O_o),
	.sel({ni11O, ni11l, ni11i, n0OOO, n0OOl, n0OOi, n0OlO}));
	defparam
		nil1O.width_data = 128,
		nil1O.width_sel = 7;
	oper_mux   nilii
	( 
	.data({{202{ni1iOli}}, 1'b1, {20{1'b0}}, 1'b1, {5{1'b0}}, 1'b1, {20{1'b0}}, 1'b1, {5{1'b0}}}),
	.o(wire_nilii_o),
	.sel({ni10l, ni11O, ni11l, ni11i, n0OOO, n0OOl, n0OOi, n0OlO}));
	defparam
		nilii.width_data = 256,
		nilii.width_sel = 8;
	oper_mux   nilil
	( 
	.data({{86{1'b0}}, 1'b1, {41{1'b0}}}),
	.o(wire_nilil_o),
	.sel({ni11O, ni11l, ni11i, n0OOO, n0OOl, n0OOi, n0OlO}));
	defparam
		nilil.width_data = 128,
		nilil.width_sel = 7;
	oper_mux   niliO
	( 
	.data({{77{1'b0}}, 1'b1, {14{1'b0}}, 1'b1, {11{1'b0}}, 1'b1, {14{1'b0}}, 1'b1, {8{1'b0}}}),
	.o(wire_niliO_o),
	.sel({ni11O, ni11l, ni11i, n0OOO, n0OOl, n0OOi, n0OlO}));
	defparam
		niliO.width_data = 128,
		niliO.width_sel = 7;
	oper_mux   nilli
	( 
	.data({{148{ni1iOli}}, {10{1'b1}}, {17{1'b0}}, 1'b1, {32{1'b0}}, 1'b1, {17{1'b0}}, 1'b1, {8{1'b0}}, 1'b1, {16{1'b0}}, 1'b1, {3{1'b0}}}),
	.o(wire_nilli_o),
	.sel({ni10l, ni11O, ni11l, ni11i, n0OOO, n0OOl, n0OOi, n0OlO}));
	defparam
		nilli.width_data = 256,
		nilli.width_sel = 8;
	oper_mux   nilll
	( 
	.data({{54{1'b0}}, 1'b1, {9{1'b0}}}),
	.o(wire_nilll_o),
	.sel({ni11O, ni11l, ni11i, n0OOO, n0OOl, n0OOi}));
	defparam
		nilll.width_data = 64,
		nilll.width_sel = 6;
	oper_mux   nillO
	( 
	.data({{81{1'b0}}, {2{1'b1}}, {45{1'b0}}}),
	.o(wire_nillO_o),
	.sel({ni11O, ni11l, ni11i, n0OOO, n0OOl, n0OOi, n0OlO}));
	defparam
		nillO.width_data = 128,
		nillO.width_sel = 7;
	oper_mux   nilOi
	( 
	.data({{56{1'b0}}, 1'b1, {71{1'b0}}}),
	.o(wire_nilOi_o),
	.sel({ni11O, ni11l, ni11i, n0OOO, n0OOl, n0OOi, n0OlO}));
	defparam
		nilOi.width_data = 128,
		nilOi.width_sel = 7;
	oper_mux   nilOl
	( 
	.data({{57{1'b0}}, 1'b1, {70{1'b0}}}),
	.o(wire_nilOl_o),
	.sel({ni11O, ni11l, ni11i, n0OOO, n0OOl, n0OOi, n0OlO}));
	defparam
		nilOl.width_data = 128,
		nilOl.width_sel = 7;
	oper_mux   nilOO
	( 
	.data({{58{1'b0}}, 1'b1, {69{1'b0}}}),
	.o(wire_nilOO_o),
	.sel({ni11O, ni11l, ni11i, n0OOO, n0OOl, n0OOi, n0OlO}));
	defparam
		nilOO.width_data = 128,
		nilOO.width_sel = 7;
	oper_mux   niO0i
	( 
	.data({{97{1'b0}}, 1'b1, {30{1'b0}}}),
	.o(wire_niO0i_o),
	.sel({ni11O, ni11l, ni11i, n0OOO, n0OOl, n0OOi, n0OlO}));
	defparam
		niO0i.width_data = 128,
		niO0i.width_sel = 7;
	oper_mux   niO0l
	( 
	.data({{98{1'b0}}, 1'b1, {29{1'b0}}}),
	.o(wire_niO0l_o),
	.sel({ni11O, ni11l, ni11i, n0OOO, n0OOl, n0OOi, n0OlO}));
	defparam
		niO0l.width_data = 128,
		niO0l.width_sel = 7;
	oper_mux   niO0O
	( 
	.data({{28{1'b0}}, {10{1'b1}}, {70{1'b0}}, {2{1'b1}}, {5{1'b0}}, {2{1'b1}}, {11{1'b0}}}),
	.o(wire_niO0O_o),
	.sel({ni11O, ni11l, ni11i, n0OOO, n0OOl, n0OOi, n0OlO}));
	defparam
		niO0O.width_data = 128,
		niO0O.width_sel = 7;
	oper_mux   niO1i
	( 
	.data({{70{1'b0}}, 1'b1, {57{1'b0}}}),
	.o(wire_niO1i_o),
	.sel({ni11O, ni11l, ni11i, n0OOO, n0OOl, n0OOi, n0OlO}));
	defparam
		niO1i.width_data = 128,
		niO1i.width_sel = 7;
	oper_mux   niO1l
	( 
	.data({{71{1'b0}}, 1'b1, {56{1'b0}}}),
	.o(wire_niO1l_o),
	.sel({ni11O, ni11l, ni11i, n0OOO, n0OOl, n0OOi, n0OlO}));
	defparam
		niO1l.width_data = 128,
		niO1l.width_sel = 7;
	oper_mux   niO1O
	( 
	.data({{26{1'b0}}, {10{1'b1}}, {45{1'b0}}, {2{1'b1}}, {5{1'b0}}, {2{1'b1}}, {38{1'b0}}}),
	.o(wire_niO1O_o),
	.sel({ni11O, ni11l, ni11i, n0OOO, n0OOl, n0OOi, n0OlO}));
	defparam
		niO1O.width_data = 128,
		niO1O.width_sel = 7;
	oper_mux   niOii
	( 
	.data({{199{ni1iOli}}, 1'b1, {54{1'b0}}, 1'b1, 1'b0}),
	.o(wire_niOii_o),
	.sel({ni10l, ni11O, ni11l, ni11i, n0OOO, n0OOl, n0OOi, n0OlO}));
	defparam
		niOii.width_data = 256,
		niOii.width_sel = 8;
	oper_mux   niOil
	( 
	.data({{157{ni1iOli}}, {10{1'b1}}, {88{1'b0}}, 1'b1}),
	.o(wire_niOil_o),
	.sel({ni10l, ni11O, ni11l, ni11i, n0OOO, n0OOl, n0OOi, n0OlO}));
	defparam
		niOil.width_data = 256,
		niOil.width_sel = 8;
	oper_mux   niOiO
	( 
	.data({{175{ni1iOli}}, 1'b1, {76{1'b0}}, 1'b1, {2{1'b0}}, 1'b1}),
	.o(wire_niOiO_o),
	.sel({ni10l, ni11O, ni11l, ni11i, n0OOO, n0OOl, n0OOi, n0OlO}));
	defparam
		niOiO.width_data = 256,
		niOiO.width_sel = 8;
	oper_mux   niOli
	( 
	.data({{175{ni1iOli}}, 1'b1, {11{1'b0}}, {2{1'b1}}, {7{1'b0}}, 1'b1, {27{1'b0}}, 1'b1, {25{1'b0}}, 1'b1, 1'b0, 1'b1, {2{1'b0}}, 1'b1}),
	.o(wire_niOli_o),
	.sel({ni10l, ni11O, ni11l, ni11i, n0OOO, n0OOl, n0OOi, n0OlO}));
	defparam
		niOli.width_data = 256,
		niOli.width_sel = 8;
	oper_mux   niOll
	( 
	.data({{124{ni1iOli}}, 1'b1, {2{1'b0}}, 1'b1, {5{1'b0}}, 1'b1, {20{1'b0}}, {10{1'b1}}, {6{1'b0}}, 1'b1, {7{1'b0}}, 1'b1, {2{1'b0}}, 1'b1, {5{1'b0}}, {2{1'b1}}, {16{1'b0}}, 1'b1, {3{1'b0}}, {2{1'b1}}, {3{1'b0}}, 1'b1, 1'b0, 1'b1, {7{1'b0}}, 1'b1, 1'b0, 1'b1, {2{1'b0}}, 1'b1, {2{1'b0}}, 1'b1, {2{1'b0}}, 1'b1, {11{1'b0}}, 1'b1, {2{1'b0}}, 1'b1, {5{1'b0}}}),
	.o(wire_niOll_o),
	.sel({ni10l, ni11O, ni11l, ni11i, n0OOO, n0OOl, n0OOi, n0OlO}));
	defparam
		niOll.width_data = 256,
		niOll.width_sel = 8;
	oper_mux   niOlO
	( 
	.data({{78{ni1iOli}}, {6{1'b1}}, {9{1'b0}}, 1'b1, 1'b0, 1'b1, {2{1'b0}}, 1'b1, {14{1'b0}}, 1'b1, {4{1'b0}}, {2{1'b1}}, 1'b0, 1'b1, {3{1'b0}}, 1'b1, {2{1'b0}}}),
	.o(wire_niOlO_o),
	.sel({ni10l, ni11O, ni11l, ni11i, n0OOO, n0OOl, n0OlO}));
	defparam
		niOlO.width_data = 128,
		niOlO.width_sel = 7;
	oper_mux   niOOi
	( 
	.data({{104{ni1iOli}}, ((ni1il0l40 ^ ni1il0l39) & ni1iOli), {3{ni1iOli}}, ((ni1il0O38 ^ ni1il0O37) & ni1iOli), {3{ni1iOli}}, ((ni1ilii36 ^ ni1ilii35) & ni1iOli), {6{ni1iOli}}, ((ni1ilil34 ^ ni1ilil33) & ni1iOli), ((ni1iliO32 ^ ni1iliO31) & ni1iOli), {77{ni1iOli}}, 1'b1, {56{1'b0}}, 1'b1}),
	.o(wire_niOOi_o),
	.sel({ni10l, ni11O, ni11l, ((ni1illi30 ^ ni1illi29) & ni11i), n0OOO, n0OOl, n0OOi, n0OlO}));
	defparam
		niOOi.width_data = 256,
		niOOi.width_sel = 8;
	oper_mux   niOOl
	( 
	.data({{4{ni1iOli}}, ((ni1illl28 ^ ni1illl27) & ni1iOli), {7{ni1iOli}}, ((ni1illO26 ^ ni1illO25) & ni1iOli), {8{ni1iOli}}, ((ni1ilOi24 ^ ni1ilOi23) & ni1iOli), {11{ni1iOli}}, ((ni1ilOl22 ^ ni1ilOl21) & ni1iOli), {8{ni1iOli}}, ((ni1ilOO20 ^ ni1ilOO19) & ni1iOli), {8{ni1iOli}}, ((ni1iO1i18 ^ ni1iO1i17) & ni1iOli), {10{ni1iOli}}, ((ni1iO1l16 ^ ni1iO1l15) & ni1iOli), {18{ni1iOli}}, ((ni1iO1O14 ^ ni1iO1O13) & ni1iOli), {7{ni1iOli}}, ((ni1iO0i12 ^ ni1iO0i11) & ni1iOli), {2{ni1iOli}}, ((ni1iO0l10 ^ ni1iO0l9) & ni1iOli), {6{ni1iOli}}, ((ni1iO0O8 ^ ni1iO0O7) & ni1iOli), ((ni1iOii6 ^ ni1iOii5) & ni1iOli), {17{ni1iOli}}, ((ni1iOil4 ^ ni1iOil3) & ni1iOli), {19{ni1iOli}}, {2{1'b1}}, {3{1'b0}}, 1'b1, {10{1'b0}}, {13{1'b1}}, {8{1'b0}}, 1'b1, {13{1'b0}}, {3{1'b1}}, {2{1'b0}}, 1'b1, {2{1'b0}}, {3{1'b1}}, {21{1'b0}}, 1'b1, {4{1'b0}}, 1'b1, {25{1'b0}}, 1'b1, {3{1'b0}}}),
	.o(wire_niOOl_o),
	.sel({ni10l, ni11O, ni11l, ni11i, n0OOO, n0OOl, n0OOi, ((ni1iOll2 ^ ni1iOll1) & n0OlO)}));
	defparam
		niOOl.width_data = 256,
		niOOl.width_sel = 8;
	oper_mux   nlO10O
	( 
	.data({{3{1'b0}}, 1'b1}),
	.o(wire_nlO10O_o),
	.sel({n110O, n110i}));
	defparam
		nlO10O.width_data = 4,
		nlO10O.width_sel = 2;
	oper_mux   nlO1ii
	( 
	.data({1'b0, 1'b1, {2{1'b0}}, 1'b1, {2{1'b0}}, 1'b1}),
	.o(wire_nlO1ii_o),
	.sel({n110O, n110l, n110i}));
	defparam
		nlO1ii.width_data = 8,
		nlO1ii.width_sel = 3;
	oper_mux   nlO1il
	( 
	.data({{2{1'b0}}, 1'b1, 1'b0, {2{1'b1}}, {2{1'b0}}}),
	.o(wire_nlO1il_o),
	.sel({n110O, n110l, n110i}));
	defparam
		nlO1il.width_data = 8,
		nlO1il.width_sel = 3;
	oper_mux   nlO1iO
	( 
	.data({1'b0, 1'b1, 1'b0, {2{1'b1}}, {3{1'b0}}}),
	.o(wire_nlO1iO_o),
	.sel({n110O, n110l, n110i}));
	defparam
		nlO1iO.width_data = 8,
		nlO1iO.width_sel = 3;
	oper_mux   nlO1li
	( 
	.data({1'b0, {2{1'b1}}, {5{1'b0}}}),
	.o(wire_nlO1li_o),
	.sel({n110O, n110l, n110i}));
	defparam
		nlO1li.width_data = 8,
		nlO1li.width_sel = 3;
	oper_mux   nlO1ll
	( 
	.data({1'b1, {7{1'b0}}}),
	.o(wire_nlO1ll_o),
	.sel({n110O, n110l, n110i}));
	defparam
		nlO1ll.width_data = 8,
		nlO1ll.width_sel = 3;
	oper_selector   ni011ii
	( 
	.data({1'b0, 1'b1, (~ nli11lO), (~ nli11OO), {14{1'b0}}}),
	.o(wire_ni011ii_o),
	.sel({1'b0, n0OOl0i, n0OOl1O, n0OOl1l, {12{1'b0}}, n0OOl1i, (~ (((n0OOl0i | n0OOl1O) | n0OOl1l) | n0OOl1i))}));
	defparam
		ni011ii.width_data = 18,
		ni011ii.width_sel = 18;
	oper_selector   ni011Ol
	( 
	.data({1'b0, 1'b1, nl0liii, nl0O01i, {14{1'b0}}}),
	.o(wire_ni011Ol_o),
	.sel({1'b0, n0OOlil, n0OOlii, n0OOl0O, {12{1'b0}}, n0OOl0l, (~ (((n0OOlil | n0OOlii) | n0OOl0O) | n0OOl0l))}));
	defparam
		ni011Ol.width_data = 18,
		ni011Ol.width_sel = 18;
	oper_selector   nii00ii
	( 
	.data({1'b0, (~ nii00li), nl00lli, {15{1'b0}}}),
	.o(wire_nii00ii_o),
	.sel({1'b0, ni1110O, ni1110l, {13{1'b0}}, ni1110i, (~ ((ni1110O | ni1110l) | ni1110i))}));
	defparam
		nii00ii.width_data = 18,
		nii00ii.width_sel = 18;
	oper_selector   nii11iO
	( 
	.data({1'b0, 1'b1, nl0liii, nl0O01i, {14{1'b0}}}),
	.o(wire_nii11iO_o),
	.sel({1'b0, n0OOOOi, n0OOOlO, n0OOOll, {12{1'b0}}, n0OOOli, (~ (((n0OOOOi | n0OOOlO) | n0OOOll) | n0OOOli))}));
	defparam
		nii11iO.width_data = 18,
		nii11iO.width_sel = 18;
	oper_selector   nii1O0O
	( 
	.data({1'b1, ni1i1il, ni1iOli}),
	.o(wire_nii1O0O_o),
	.sel({(~ n0Oll), n0Oll, 1'b0}));
	defparam
		nii1O0O.width_data = 3,
		nii1O0O.width_sel = 3;
	oper_selector   nil10iO
	( 
	.data({1'b0, (((~ nil10lO) & nl1OOll) & nl1OOOl), ((nl1i0OO | nl1i0Oi) & (~ nil10lO)), (~ nil10lO), nl00O0i, {13{1'b0}}}),
	.o(wire_nil10iO_o),
	.sel({1'b0, ni1100O, ni1100l, ni1100i, ni1101O, {11{1'b0}}, ni1101l, (~ ni1101i)}));
	defparam
		nil10iO.width_data = 18,
		nil10iO.width_sel = 18;
	oper_selector   nilOill
	( 
	.data({1'b0, (~ nilOiOl), (((nl1OOll & nl0l11l) & nl1OOOl) & (~ nilOiOl)), ((nl1i0OO | nl1i0Oi) & (~ nilOiOl)), (nl1i0OO | nl1i0Oi), {13{1'b0}}}),
	.o(wire_nilOill_o),
	.sel({1'b0, ni11i0O, ni11i0l, ni11i0i, ni11i1O, {11{1'b0}}, ni11i1l, (~ ni11i1i)}));
	defparam
		nilOill.width_data = 18,
		nilOill.width_sel = 18;
	oper_selector   niO0i1l
	( 
	.data({1'b1, (~ nl0lili), (((nl0l1ll & nl0li0i) | (~ nl0li0i)) & (~ nl0lili)), {15{1'b0}}}),
	.o(wire_niO0i1l_o),
	.sel({ni11l0i, ni11l1O, ni11l1l, {13{1'b0}}, ni11l1i, (~ (((ni11l0i | ni11l1O) | ni11l1l) | ni11l1i))}));
	defparam
		niO0i1l.width_data = 18,
		niO0i1l.width_sel = 18;
	oper_selector   niO0ili
	( 
	.data({1'b0, 1'b1, nl0lili, ni1iiOi, ni1iilO, {13{1'b0}}}),
	.o(wire_niO0ili_o),
	.sel({1'b0, ni11lli, ni11liO, ni11lil, ni11lii, {11{1'b0}}, ni11l0O, (~ ni11l0l)}));
	defparam
		niO0ili.width_data = 18,
		niO0ili.width_sel = 18;
	oper_selector   niO0O0O
	( 
	.data({nii11lO, nli0O1l, ni1iOli}),
	.o(wire_niO0O0O_o),
	.sel({(~ n11li), n11li, 1'b0}));
	defparam
		niO0O0O.width_data = 3,
		niO0O0O.width_sel = 3;
	oper_selector   niO0Oii
	( 
	.data({nii11Oi, nli0O1O, ni1iOli}),
	.o(wire_niO0Oii_o),
	.sel({(~ n11li), n11li, 1'b0}));
	defparam
		niO0Oii.width_data = 3,
		niO0Oii.width_sel = 3;
	oper_selector   niO0Oil
	( 
	.data({nii11Ol, nli0O0i, ni1iOli}),
	.o(wire_niO0Oil_o),
	.sel({(~ n11li), n11li, 1'b0}));
	defparam
		niO0Oil.width_data = 3,
		niO0Oil.width_sel = 3;
	oper_selector   niO0OiO
	( 
	.data({nii11OO, nli0O0l, ni1iOli}),
	.o(wire_niO0OiO_o),
	.sel({(~ n11li), n11li, 1'b0}));
	defparam
		niO0OiO.width_data = 3,
		niO0OiO.width_sel = 3;
	oper_selector   niO0Oli
	( 
	.data({nii101i, nli0O0O, ni1iOli}),
	.o(wire_niO0Oli_o),
	.sel({(~ n11li), n11li, 1'b0}));
	defparam
		niO0Oli.width_data = 3,
		niO0Oli.width_sel = 3;
	oper_selector   niO0Oll
	( 
	.data({nii101l, nli0Oii, ni1iOli}),
	.o(wire_niO0Oll_o),
	.sel({(~ n11li), n11li, 1'b0}));
	defparam
		niO0Oll.width_data = 3,
		niO0Oll.width_sel = 3;
	oper_selector   niO0OlO
	( 
	.data({nii101O, nli0Oil, ni1iOli}),
	.o(wire_niO0OlO_o),
	.sel({(~ n11li), n11li, 1'b0}));
	defparam
		niO0OlO.width_data = 3,
		niO0OlO.width_sel = 3;
	oper_selector   niO0OOi
	( 
	.data({nii100i, nli0OiO, ni1iOli}),
	.o(wire_niO0OOi_o),
	.sel({(~ n11li), n11li, 1'b0}));
	defparam
		niO0OOi.width_data = 3,
		niO0OOi.width_sel = 3;
	oper_selector   niO0OOl
	( 
	.data({nii100l, nli0Oli, ni1iOli}),
	.o(wire_niO0OOl_o),
	.sel({(~ n11li), n11li, 1'b0}));
	defparam
		niO0OOl.width_data = 3,
		niO0OOl.width_sel = 3;
	oper_selector   niO0OOO
	( 
	.data({nii100O, nli0Oll, ni1iOli}),
	.o(wire_niO0OOO_o),
	.sel({(~ n11li), n11li, 1'b0}));
	defparam
		niO0OOO.width_data = 3,
		niO0OOO.width_sel = 3;
	oper_selector   niOi00O
	( 
	.data({1'b0, 1'b1, nl0lili, ni1iiOi, ni1iilO, {13{1'b0}}}),
	.o(wire_niOi00O_o),
	.sel({1'b0, ni11O1i, ni11lOO, ni11lOl, ni11lOi, {11{1'b0}}, ni11llO, (~ ni11lll)}));
	defparam
		niOi00O.width_data = 18,
		niOi00O.width_sel = 18;
	oper_selector   niOi0Oi
	( 
	.data({1'b1, nl0lili, nii1iii, {15{1'b0}}}),
	.o(wire_niOi0Oi_o),
	.sel({ni11O0l, ni11O0i, ni11O1O, {13{1'b0}}, ni11O1l, (~ (((ni11O0l | ni11O0i) | ni11O1O) | ni11O1l))}));
	defparam
		niOi0Oi.width_data = 18,
		niOi0Oi.width_sel = 18;
	oper_selector   niOi10i
	( 
	.data({nii10li, nli0OOO, ni1iOli}),
	.o(wire_niOi10i_o),
	.sel({(~ n11li), n11li, 1'b0}));
	defparam
		niOi10i.width_data = 3,
		niOi10i.width_sel = 3;
	oper_selector   niOi10l
	( 
	.data({nii10ll, nlii11i, ni1iOli}),
	.o(wire_niOi10l_o),
	.sel({(~ n11li), n11li, 1'b0}));
	defparam
		niOi10l.width_data = 3,
		niOi10l.width_sel = 3;
	oper_selector   niOi10O
	( 
	.data({nii10lO, nlii11l, ni1iOli}),
	.o(wire_niOi10O_o),
	.sel({(~ n11li), n11li, 1'b0}));
	defparam
		niOi10O.width_data = 3,
		niOi10O.width_sel = 3;
	oper_selector   niOi11i
	( 
	.data({nii10ii, nli0OlO, ni1iOli}),
	.o(wire_niOi11i_o),
	.sel({(~ n11li), n11li, 1'b0}));
	defparam
		niOi11i.width_data = 3,
		niOi11i.width_sel = 3;
	oper_selector   niOi11l
	( 
	.data({nii10il, nli0OOi, ni1iOli}),
	.o(wire_niOi11l_o),
	.sel({(~ n11li), n11li, 1'b0}));
	defparam
		niOi11l.width_data = 3,
		niOi11l.width_sel = 3;
	oper_selector   niOi11O
	( 
	.data({nii10iO, nli0OOl, ni1iOli}),
	.o(wire_niOi11O_o),
	.sel({(~ n11li), n11li, 1'b0}));
	defparam
		niOi11O.width_data = 3,
		niOi11O.width_sel = 3;
	oper_selector   niOi1ii
	( 
	.data({nii10Oi, nlii11O, ni1iOli}),
	.o(wire_niOi1ii_o),
	.sel({(~ n11li), n11li, 1'b0}));
	defparam
		niOi1ii.width_data = 3,
		niOi1ii.width_sel = 3;
	oper_selector   niOi1il
	( 
	.data({nii10Ol, nlii10i, ni1iOli}),
	.o(wire_niOi1il_o),
	.sel({(~ n11li), n11li, 1'b0}));
	defparam
		niOi1il.width_data = 3,
		niOi1il.width_sel = 3;
	oper_selector   niOi1iO
	( 
	.data({nii10OO, nlii10l, ni1iOli}),
	.o(wire_niOi1iO_o),
	.sel({(~ n11li), n11li, 1'b0}));
	defparam
		niOi1iO.width_data = 3,
		niOi1iO.width_sel = 3;
	oper_selector   niOi1li
	( 
	.data({nii1i1i, nlii10O, ni1iOli}),
	.o(wire_niOi1li_o),
	.sel({(~ n11li), n11li, 1'b0}));
	defparam
		niOi1li.width_data = 3,
		niOi1li.width_sel = 3;
	oper_selector   niOi1ll
	( 
	.data({nii1i1l, nlii1ii, ni1iOli}),
	.o(wire_niOi1ll_o),
	.sel({(~ n11li), n11li, 1'b0}));
	defparam
		niOi1ll.width_data = 3,
		niOi1ll.width_sel = 3;
	oper_selector   niOi1lO
	( 
	.data({nii1i1O, nlii1il, ni1iOli}),
	.o(wire_niOi1lO_o),
	.sel({(~ n11li), n11li, 1'b0}));
	defparam
		niOi1lO.width_data = 3,
		niOi1lO.width_sel = 3;
	oper_selector   niOi1Oi
	( 
	.data({nii1i0i, nlii1iO, ni1iOli}),
	.o(wire_niOi1Oi_o),
	.sel({(~ n11li), n11li, 1'b0}));
	defparam
		niOi1Oi.width_data = 3,
		niOi1Oi.width_sel = 3;
	oper_selector   niOi1Ol
	( 
	.data({nii1i0l, nlii1ll, ni1iOli}),
	.o(wire_niOi1Ol_o),
	.sel({(~ n11li), n11li, 1'b0}));
	defparam
		niOi1Ol.width_data = 3,
		niOi1Ol.width_sel = 3;
	oper_selector   niOll0O
	( 
	.data({1'b0, nl10l0O, ni1iOli}),
	.o(wire_niOll0O_o),
	.sel({(~ n0Oll), n0Oll, 1'b0}));
	defparam
		niOll0O.width_data = 3,
		niOll0O.width_sel = 3;
	oper_selector   niOllii
	( 
	.data({1'b0, nl10lii, ni1iOli}),
	.o(wire_niOllii_o),
	.sel({(~ n0Oll), n0Oll, 1'b0}));
	defparam
		niOllii.width_data = 3,
		niOllii.width_sel = 3;
	oper_selector   niOllil
	( 
	.data({1'b0, nl10lil, ni1iOli}),
	.o(wire_niOllil_o),
	.sel({(~ n0Oll), n0Oll, 1'b0}));
	defparam
		niOllil.width_data = 3,
		niOllil.width_sel = 3;
	oper_selector   niOlliO
	( 
	.data({1'b0, nl10liO, ni1iOli}),
	.o(wire_niOlliO_o),
	.sel({(~ n0Oll), n0Oll, 1'b0}));
	defparam
		niOlliO.width_data = 3,
		niOlliO.width_sel = 3;
	oper_selector   niOllli
	( 
	.data({1'b0, nl10lli, ni1iOli}),
	.o(wire_niOllli_o),
	.sel({(~ n0Oll), n0Oll, 1'b0}));
	defparam
		niOllli.width_data = 3,
		niOllli.width_sel = 3;
	oper_selector   niOllll
	( 
	.data({1'b0, nl10lll, ni1iOli}),
	.o(wire_niOllll_o),
	.sel({(~ n0Oll), n0Oll, 1'b0}));
	defparam
		niOllll.width_data = 3,
		niOllll.width_sel = 3;
	oper_selector   niOlllO
	( 
	.data({1'b0, nl10llO, ni1iOli}),
	.o(wire_niOlllO_o),
	.sel({(~ n0Oll), n0Oll, 1'b0}));
	defparam
		niOlllO.width_data = 3,
		niOlllO.width_sel = 3;
	oper_selector   niOllOi
	( 
	.data({1'b0, nl10lOi, ni1iOli}),
	.o(wire_niOllOi_o),
	.sel({(~ n0Oll), n0Oll, 1'b0}));
	defparam
		niOllOi.width_data = 3,
		niOllOi.width_sel = 3;
	oper_selector   niOllOl
	( 
	.data({1'b0, nl10lOO, ni1iOli}),
	.o(wire_niOllOl_o),
	.sel({(~ n0Oll), n0Oll, 1'b0}));
	defparam
		niOllOl.width_data = 3,
		niOllOl.width_sel = 3;
	oper_selector   niOllOO
	( 
	.data({1'b0, nl10O1l, ni1iOli}),
	.o(wire_niOllOO_o),
	.sel({(~ n0Oll), n0Oll, 1'b0}));
	defparam
		niOllOO.width_data = 3,
		niOllOO.width_sel = 3;
	oper_selector   niOlOOl
	( 
	.data({1'b0, nl0i10l, ni1iOli}),
	.o(wire_niOlOOl_o),
	.sel({(~ n0lli), n0lli, 1'b0}));
	defparam
		niOlOOl.width_data = 3,
		niOlOOl.width_sel = 3;
	oper_selector   niOO0iO
	( 
	.data({1'b0, nl0i10l, ni1iOli}),
	.o(wire_niOO0iO_o),
	.sel({(~ n0liO), n0liO, 1'b0}));
	defparam
		niOO0iO.width_data = 3,
		niOO0iO.width_sel = 3;
	oper_selector   niOOlOO
	( 
	.data({1'b0, nii0i1i, ni1iOli}),
	.o(wire_niOOlOO_o),
	.sel({(~ n0OiO), n0OiO, 1'b0}));
	defparam
		niOOlOO.width_data = 3,
		niOOlOO.width_sel = 3;
	oper_selector   niOOO0i
	( 
	.data({1'b0, nii0i0l, ni1iOli}),
	.o(wire_niOOO0i_o),
	.sel({(~ n0OiO), n0OiO, 1'b0}));
	defparam
		niOOO0i.width_data = 3,
		niOOO0i.width_sel = 3;
	oper_selector   niOOO0l
	( 
	.data({1'b0, nii0i0O, ni1iOli}),
	.o(wire_niOOO0l_o),
	.sel({(~ n0OiO), n0OiO, 1'b0}));
	defparam
		niOOO0l.width_data = 3,
		niOOO0l.width_sel = 3;
	oper_selector   niOOO0O
	( 
	.data({1'b0, nii0iii, ni1iOli}),
	.o(wire_niOOO0O_o),
	.sel({(~ n0OiO), n0OiO, 1'b0}));
	defparam
		niOOO0O.width_data = 3,
		niOOO0O.width_sel = 3;
	oper_selector   niOOO1i
	( 
	.data({1'b0, nii0i1l, ni1iOli}),
	.o(wire_niOOO1i_o),
	.sel({(~ n0OiO), n0OiO, 1'b0}));
	defparam
		niOOO1i.width_data = 3,
		niOOO1i.width_sel = 3;
	oper_selector   niOOO1l
	( 
	.data({1'b0, nii0i1O, ni1iOli}),
	.o(wire_niOOO1l_o),
	.sel({(~ n0OiO), n0OiO, 1'b0}));
	defparam
		niOOO1l.width_data = 3,
		niOOO1l.width_sel = 3;
	oper_selector   niOOO1O
	( 
	.data({1'b0, nii0i0i, ni1iOli}),
	.o(wire_niOOO1O_o),
	.sel({(~ n0OiO), n0OiO, 1'b0}));
	defparam
		niOOO1O.width_data = 3,
		niOOO1O.width_sel = 3;
	oper_selector   niOOOii
	( 
	.data({1'b0, nii0iil, ni1iOli}),
	.o(wire_niOOOii_o),
	.sel({(~ n0OiO), n0OiO, 1'b0}));
	defparam
		niOOOii.width_data = 3,
		niOOOii.width_sel = 3;
	oper_selector   niOOOil
	( 
	.data({1'b0, nii0iiO, ni1iOli}),
	.o(wire_niOOOil_o),
	.sel({(~ n0OiO), n0OiO, 1'b0}));
	defparam
		niOOOil.width_data = 3,
		niOOOil.width_sel = 3;
	oper_selector   niOOOiO
	( 
	.data({1'b0, nii0ili, ni1iOli}),
	.o(wire_niOOOiO_o),
	.sel({(~ n0OiO), n0OiO, 1'b0}));
	defparam
		niOOOiO.width_data = 3,
		niOOOiO.width_sel = 3;
	oper_selector   niOOOli
	( 
	.data({1'b0, nii0ill, ni1iOli}),
	.o(wire_niOOOli_o),
	.sel({(~ n0OiO), n0OiO, 1'b0}));
	defparam
		niOOOli.width_data = 3,
		niOOOli.width_sel = 3;
	oper_selector   niOOOll
	( 
	.data({1'b0, nii0ilO, ni1iOli}),
	.o(wire_niOOOll_o),
	.sel({(~ n0OiO), n0OiO, 1'b0}));
	defparam
		niOOOll.width_data = 3,
		niOOOll.width_sel = 3;
	oper_selector   niOOOlO
	( 
	.data({1'b0, nii0iOi, ni1iOli}),
	.o(wire_niOOOlO_o),
	.sel({(~ n0OiO), n0OiO, 1'b0}));
	defparam
		niOOOlO.width_data = 3,
		niOOOlO.width_sel = 3;
	oper_selector   niOOOOi
	( 
	.data({1'b0, nii0iOl, ni1iOli}),
	.o(wire_niOOOOi_o),
	.sel({(~ n0OiO), n0OiO, 1'b0}));
	defparam
		niOOOOi.width_data = 3,
		niOOOOi.width_sel = 3;
	oper_selector   niOOOOl
	( 
	.data({1'b0, nii0iOO, ni1iOli}),
	.o(wire_niOOOOl_o),
	.sel({(~ n0OiO), n0OiO, 1'b0}));
	defparam
		niOOOOl.width_data = 3,
		niOOOOl.width_sel = 3;
	oper_selector   niOOOOO
	( 
	.data({1'b0, nii0l1i, ni1iOli}),
	.o(wire_niOOOOO_o),
	.sel({(~ n0OiO), n0OiO, 1'b0}));
	defparam
		niOOOOO.width_data = 3,
		niOOOOO.width_sel = 3;
	oper_selector   nl000iO
	( 
	.data({1'b0, niOlOlO, ni1iOli}),
	.o(wire_nl000iO_o),
	.sel({(~ n0Oll), n0Oll, 1'b0}));
	defparam
		nl000iO.width_data = 3,
		nl000iO.width_sel = 3;
	oper_selector   nl000li
	( 
	.data({1'b0, niOlO1l, ni1iOli}),
	.o(wire_nl000li_o),
	.sel({(~ n0Oll), n0Oll, 1'b0}));
	defparam
		nl000li.width_data = 3,
		nl000li.width_sel = 3;
	oper_selector   nl000ll
	( 
	.data({1'b0, niOlO1O, ni1iOli}),
	.o(wire_nl000ll_o),
	.sel({(~ n0Oll), n0Oll, 1'b0}));
	defparam
		nl000ll.width_data = 3,
		nl000ll.width_sel = 3;
	oper_selector   nl000lO
	( 
	.data({1'b0, niOlO0i, ni1iOli}),
	.o(wire_nl000lO_o),
	.sel({(~ n0Oll), n0Oll, 1'b0}));
	defparam
		nl000lO.width_data = 3,
		nl000lO.width_sel = 3;
	oper_selector   nl000Oi
	( 
	.data({1'b0, niOlO0l, ni1iOli}),
	.o(wire_nl000Oi_o),
	.sel({(~ n0Oll), n0Oll, 1'b0}));
	defparam
		nl000Oi.width_data = 3,
		nl000Oi.width_sel = 3;
	oper_selector   nl000Ol
	( 
	.data({1'b0, niOlO0O, ni1iOli}),
	.o(wire_nl000Ol_o),
	.sel({(~ n0Oll), n0Oll, 1'b0}));
	defparam
		nl000Ol.width_data = 3,
		nl000Ol.width_sel = 3;
	oper_selector   nl000OO
	( 
	.data({1'b0, niOlOii, ni1iOli}),
	.o(wire_nl000OO_o),
	.sel({(~ n0Oll), n0Oll, 1'b0}));
	defparam
		nl000OO.width_data = 3,
		nl000OO.width_sel = 3;
	oper_selector   nl0010O
	( 
	.data({1'b0, 1'b1, nl0lili, nl0lOOi, (~ nl0lili), (~ nl0l1Oi), nii1iii, (~ nii1iii), nl0li1i, {9{1'b0}}}),
	.o(wire_nl0010O_o),
	.sel({1'b0, ni10O1i, ni10lOO, ni10lOl, ni10lOi, ni10llO, ni10lll, ni10lli, ni10liO, {7{1'b0}}, ni10lil, (~ ni10lii)}));
	defparam
		nl0010O.width_data = 18,
		nl0010O.width_sel = 18;
	oper_selector   nl00i1i
	( 
	.data({1'b0, niOlOil, ni1iOli}),
	.o(wire_nl00i1i_o),
	.sel({(~ n0Oll), n0Oll, 1'b0}));
	defparam
		nl00i1i.width_data = 3,
		nl00i1i.width_sel = 3;
	oper_selector   nl00i1l
	( 
	.data({1'b0, niOlOiO, ni1iOli}),
	.o(wire_nl00i1l_o),
	.sel({(~ n0Oll), n0Oll, 1'b0}));
	defparam
		nl00i1l.width_data = 3,
		nl00i1l.width_sel = 3;
	oper_selector   nl00i1O
	( 
	.data({1'b0, niOlOli, ni1iOli}),
	.o(wire_nl00i1O_o),
	.sel({(~ n0Oll), n0Oll, 1'b0}));
	defparam
		nl00i1O.width_data = 3,
		nl00i1O.width_sel = 3;
	oper_selector   nl010ll
	( 
	.data({nii11lO, nlii01i, ni1iOli}),
	.o(wire_nl010ll_o),
	.sel({(~ n111l), n111l, 1'b0}));
	defparam
		nl010ll.width_data = 3,
		nl010ll.width_sel = 3;
	oper_selector   nl010lO
	( 
	.data({nii11Oi, nlii01l, ni1iOli}),
	.o(wire_nl010lO_o),
	.sel({(~ n111l), n111l, 1'b0}));
	defparam
		nl010lO.width_data = 3,
		nl010lO.width_sel = 3;
	oper_selector   nl010Oi
	( 
	.data({nii11Ol, nlii01O, ni1iOli}),
	.o(wire_nl010Oi_o),
	.sel({(~ n111l), n111l, 1'b0}));
	defparam
		nl010Oi.width_data = 3,
		nl010Oi.width_sel = 3;
	oper_selector   nl010Ol
	( 
	.data({nii11OO, nlii00l, ni1iOli}),
	.o(wire_nl010Ol_o),
	.sel({(~ n111l), n111l, 1'b0}));
	defparam
		nl010Ol.width_data = 3,
		nl010Ol.width_sel = 3;
	oper_selector   nl0111l
	( 
	.data({nlii01i, nlii0Oi, ni1iOli}),
	.o(wire_nl0111l_o),
	.sel({(~ n10li), n10li, 1'b0}));
	defparam
		nl0111l.width_data = 3,
		nl0111l.width_sel = 3;
	oper_selector   nl0111O
	( 
	.data({nlii01l, nlii0Ol, ni1iOli}),
	.o(wire_nl0111O_o),
	.sel({(~ n10li), n10li, 1'b0}));
	defparam
		nl0111O.width_data = 3,
		nl0111O.width_sel = 3;
	oper_selector   nl011lO
	( 
	.data({nii11lO, nlii0Oi, ni1iOli}),
	.o(wire_nl011lO_o),
	.sel({(~ n10li), n10li, 1'b0}));
	defparam
		nl011lO.width_data = 3,
		nl011lO.width_sel = 3;
	oper_selector   nl011Oi
	( 
	.data({nii11Oi, nlii0Ol, ni1iOli}),
	.o(wire_nl011Oi_o),
	.sel({(~ n10li), n10li, 1'b0}));
	defparam
		nl011Oi.width_data = 3,
		nl011Oi.width_sel = 3;
	oper_selector   nl011Ol
	( 
	.data({nii11Ol, nlii0OO, ni1iOli}),
	.o(wire_nl011Ol_o),
	.sel({(~ n10li), n10li, 1'b0}));
	defparam
		nl011Ol.width_data = 3,
		nl011Ol.width_sel = 3;
	oper_selector   nl011OO
	( 
	.data({nii11OO, nliii1l, ni1iOli}),
	.o(wire_nl011OO_o),
	.sel({(~ n10li), n10li, 1'b0}));
	defparam
		nl011OO.width_data = 3,
		nl011OO.width_sel = 3;
	oper_selector   nl01lii
	( 
	.data({1'b0, 1'b1, nl0i0ll, (~ ni10Oll), (~ ni10OlO), (~ wire_niOl0il_q_a[0]), (~ ni10OOi), (~ ((~ nii00li) & (~ ni10Oll))), nilOiOl, (~ ((~ nii00li) & wire_nl0O00O_o[9])), (~ wire_nl0O0ii_o[11]), ((~ nii00li) & wire_nl0O00O_o[9]), (~ nl0l0il), (~ ((~ nil10lO) & (~ ni10OlO))), nl0l0il, {3{1'b0}}}),
	.o(wire_nl01lii_o),
	.sel({1'b0, ni10iOl, ni10iOi, ni10ilO, ni10ill, ni10ili, ni10iiO, ni10iil, ni10iii, ni10i0O, ni10i0l, ni10i0i, ni10i1O, ni10i1l, ni10i1i, 1'b0, ni100OO, (~ ni100Ol)}));
	defparam
		nl01lii.width_data = 18,
		nl01lii.width_sel = 18;
	oper_selector   nl01O1i
	( 
	.data({1'b0, wire_nl0O0ii_o[11], ((~ nii00li) & (~ ni10Oll)), (~ nilOiOl), (~ nl0i0Oi), ((~ nil10lO) & (~ ni10OlO)), {12{1'b0}}}),
	.o(wire_nl01O1i_o),
	.sel({1'b0, ni10l0O, ni10l0l, ni10l0i, ni10l1O, ni10l1l, {10{1'b0}}, ni10l1i, (~ ni10iOO)}));
	defparam
		nl01O1i.width_data = 18,
		nl01O1i.width_sel = 18;
	oper_selector   nl01Oli
	( 
	.data({1'b0, (~ nl0lOOi), ni1iOli}),
	.o(wire_nl01Oli_o),
	.sel({(~ n10Ol), n10Ol, 1'b0}));
	defparam
		nl01Oli.width_data = 3,
		nl01Oli.width_sel = 3;
	oper_selector   nl0l00l
	( 
	.data({1'b0, 1'b1, ni1iOli}),
	.o(wire_nl0l00l_o),
	.sel({(~ n11li), n11li, 1'b0}));
	defparam
		nl0l00l.width_data = 3,
		nl0l00l.width_sel = 3;
	oper_selector   nl0l0li
	( 
	.data({(nl0li0i | nlii1Ol), nl0l0il, ni1iOli}),
	.o(wire_nl0l0li_o),
	.sel({(~ n11ll), n11ll, 1'b0}));
	defparam
		nl0l0li.width_data = 3,
		nl0l0li.width_sel = 3;
	oper_selector   nl0llii
	( 
	.data({nl00i0l, nl0lOOO, ni1iOli}),
	.o(wire_nl0llii_o),
	.sel({(~ n11li), n11li, 1'b0}));
	defparam
		nl0llii.width_data = 3,
		nl0llii.width_sel = 3;
	oper_selector   nl0llil
	( 
	.data({nl00i0O, nl0lO0i, ni1iOli}),
	.o(wire_nl0llil_o),
	.sel({(~ n11li), n11li, 1'b0}));
	defparam
		nl0llil.width_data = 3,
		nl0llil.width_sel = 3;
	oper_selector   nl0lliO
	( 
	.data({nl00iii, nl0lO0l, ni1iOli}),
	.o(wire_nl0lliO_o),
	.sel({(~ n11li), n11li, 1'b0}));
	defparam
		nl0lliO.width_data = 3,
		nl0lliO.width_sel = 3;
	oper_selector   nl0llli
	( 
	.data({nl00iil, nl0lO0O, ni1iOli}),
	.o(wire_nl0llli_o),
	.sel({(~ n11li), n11li, 1'b0}));
	defparam
		nl0llli.width_data = 3,
		nl0llli.width_sel = 3;
	oper_selector   nl0llll
	( 
	.data({nl00iiO, nl0lOii, ni1iOli}),
	.o(wire_nl0llll_o),
	.sel({(~ n11li), n11li, 1'b0}));
	defparam
		nl0llll.width_data = 3,
		nl0llll.width_sel = 3;
	oper_selector   nl0lllO
	( 
	.data({nl00ili, nl0lOil, ni1iOli}),
	.o(wire_nl0lllO_o),
	.sel({(~ n11li), n11li, 1'b0}));
	defparam
		nl0lllO.width_data = 3,
		nl0lllO.width_sel = 3;
	oper_selector   nl0llOi
	( 
	.data({nl00ill, nl0lOiO, ni1iOli}),
	.o(wire_nl0llOi_o),
	.sel({(~ n11li), n11li, 1'b0}));
	defparam
		nl0llOi.width_data = 3,
		nl0llOi.width_sel = 3;
	oper_selector   nl0llOl
	( 
	.data({nl00ilO, nl0lOli, ni1iOli}),
	.o(wire_nl0llOl_o),
	.sel({(~ n11li), n11li, 1'b0}));
	defparam
		nl0llOl.width_data = 3,
		nl0llOl.width_sel = 3;
	oper_selector   nl0llOO
	( 
	.data({nl00iOi, nl0lOll, ni1iOli}),
	.o(wire_nl0llOO_o),
	.sel({(~ n11li), n11li, 1'b0}));
	defparam
		nl0llOO.width_data = 3,
		nl0llOO.width_sel = 3;
	oper_selector   nl0lO1i
	( 
	.data({nl00iOO, nl0lOlO, ni1iOli}),
	.o(wire_nl0lO1i_o),
	.sel({(~ n11li), n11li, 1'b0}));
	defparam
		nl0lO1i.width_data = 3,
		nl0lO1i.width_sel = 3;
	oper_selector   nl0lO1l
	( 
	.data({1'b0, nl0lOOi, ni1iOli}),
	.o(wire_nl0lO1l_o),
	.sel({(~ n11li), n11li, 1'b0}));
	defparam
		nl0lO1l.width_data = 3,
		nl0lO1l.width_sel = 3;
	oper_selector   nl1000O
	( 
	.data({1'b1, (~ nli11OO), nl00O0i, {15{1'b0}}}),
	.o(wire_nl1000O_o),
	.sel({ni101li, ni101iO, ni101il, {13{1'b0}}, ni101ii, (~ (((ni101li | ni101iO) | ni101il) | ni101ii))}));
	defparam
		nl1000O.width_data = 18,
		nl1000O.width_sel = 18;
	oper_selector   nl1010i
	( 
	.data({1'b0, nil1iOO, ni1iOli}),
	.o(wire_nl1010i_o),
	.sel({(~ n0Oil), n0Oil, 1'b0}));
	defparam
		nl1010i.width_data = 3,
		nl1010i.width_sel = 3;
	oper_selector   nl1010l
	( 
	.data({1'b0, nil1l1i, ni1iOli}),
	.o(wire_nl1010l_o),
	.sel({(~ n0Oil), n0Oil, 1'b0}));
	defparam
		nl1010l.width_data = 3,
		nl1010l.width_sel = 3;
	oper_selector   nl1010O
	( 
	.data({1'b0, nil1l1l, ni1iOli}),
	.o(wire_nl1010O_o),
	.sel({(~ n0Oil), n0Oil, 1'b0}));
	defparam
		nl1010O.width_data = 3,
		nl1010O.width_sel = 3;
	oper_selector   nl1011i
	( 
	.data({1'b0, nil1ilO, ni1iOli}),
	.o(wire_nl1011i_o),
	.sel({(~ n0Oil), n0Oil, 1'b0}));
	defparam
		nl1011i.width_data = 3,
		nl1011i.width_sel = 3;
	oper_selector   nl1011l
	( 
	.data({1'b0, nil1iOi, ni1iOli}),
	.o(wire_nl1011l_o),
	.sel({(~ n0Oil), n0Oil, 1'b0}));
	defparam
		nl1011l.width_data = 3,
		nl1011l.width_sel = 3;
	oper_selector   nl1011O
	( 
	.data({1'b0, nil1iOl, ni1iOli}),
	.o(wire_nl1011O_o),
	.sel({(~ n0Oil), n0Oil, 1'b0}));
	defparam
		nl1011O.width_data = 3,
		nl1011O.width_sel = 3;
	oper_selector   nl101ii
	( 
	.data({1'b0, nil1l1O, ni1iOli}),
	.o(wire_nl101ii_o),
	.sel({(~ n0Oil), n0Oil, 1'b0}));
	defparam
		nl101ii.width_data = 3,
		nl101ii.width_sel = 3;
	oper_selector   nl101il
	( 
	.data({1'b0, nil1l0i, ni1iOli}),
	.o(wire_nl101il_o),
	.sel({(~ n0Oil), n0Oil, 1'b0}));
	defparam
		nl101il.width_data = 3,
		nl101il.width_sel = 3;
	oper_selector   nl101iO
	( 
	.data({1'b0, nil1l0l, ni1iOli}),
	.o(wire_nl101iO_o),
	.sel({(~ n0Oil), n0Oil, 1'b0}));
	defparam
		nl101iO.width_data = 3,
		nl101iO.width_sel = 3;
	oper_selector   nl101li
	( 
	.data({1'b0, nil1l0O, ni1iOli}),
	.o(wire_nl101li_o),
	.sel({(~ n0Oil), n0Oil, 1'b0}));
	defparam
		nl101li.width_data = 3,
		nl101li.width_sel = 3;
	oper_selector   nl101ll
	( 
	.data({1'b0, nil1lii, ni1iOli}),
	.o(wire_nl101ll_o),
	.sel({(~ n0Oil), n0Oil, 1'b0}));
	defparam
		nl101ll.width_data = 3,
		nl101ll.width_sel = 3;
	oper_selector   nl101lO
	( 
	.data({1'b0, nil1lil, ni1iOli}),
	.o(wire_nl101lO_o),
	.sel({(~ n0Oil), n0Oil, 1'b0}));
	defparam
		nl101lO.width_data = 3,
		nl101lO.width_sel = 3;
	oper_selector   nl101Oi
	( 
	.data({1'b0, nil1liO, ni1iOli}),
	.o(wire_nl101Oi_o),
	.sel({(~ n0Oil), n0Oil, 1'b0}));
	defparam
		nl101Oi.width_data = 3,
		nl101Oi.width_sel = 3;
	oper_selector   nl101Ol
	( 
	.data({1'b0, nil1lli, ni1iOli}),
	.o(wire_nl101Ol_o),
	.sel({(~ n0Oil), n0Oil, 1'b0}));
	defparam
		nl101Ol.width_data = 3,
		nl101Ol.width_sel = 3;
	oper_selector   nl101OO
	( 
	.data({1'b0, nil1llO, ni1iOli}),
	.o(wire_nl101OO_o),
	.sel({(~ n0Oil), n0Oil, 1'b0}));
	defparam
		nl101OO.width_data = 3,
		nl101OO.width_sel = 3;
	oper_selector   nl1110i
	( 
	.data({1'b0, nii0l0l, ni1iOli}),
	.o(wire_nl1110i_o),
	.sel({(~ n0OiO), n0OiO, 1'b0}));
	defparam
		nl1110i.width_data = 3,
		nl1110i.width_sel = 3;
	oper_selector   nl1110l
	( 
	.data({1'b0, nii0l0O, ni1iOli}),
	.o(wire_nl1110l_o),
	.sel({(~ n0OiO), n0OiO, 1'b0}));
	defparam
		nl1110l.width_data = 3,
		nl1110l.width_sel = 3;
	oper_selector   nl1110O
	( 
	.data({1'b0, nii0lii, ni1iOli}),
	.o(wire_nl1110O_o),
	.sel({(~ n0OiO), n0OiO, 1'b0}));
	defparam
		nl1110O.width_data = 3,
		nl1110O.width_sel = 3;
	oper_selector   nl1111i
	( 
	.data({1'b0, nii0l1l, ni1iOli}),
	.o(wire_nl1111i_o),
	.sel({(~ n0OiO), n0OiO, 1'b0}));
	defparam
		nl1111i.width_data = 3,
		nl1111i.width_sel = 3;
	oper_selector   nl1111l
	( 
	.data({1'b0, nii0l1O, ni1iOli}),
	.o(wire_nl1111l_o),
	.sel({(~ n0OiO), n0OiO, 1'b0}));
	defparam
		nl1111l.width_data = 3,
		nl1111l.width_sel = 3;
	oper_selector   nl1111O
	( 
	.data({1'b0, nii0l0i, ni1iOli}),
	.o(wire_nl1111O_o),
	.sel({(~ n0OiO), n0OiO, 1'b0}));
	defparam
		nl1111O.width_data = 3,
		nl1111O.width_sel = 3;
	oper_selector   nl111ii
	( 
	.data({1'b0, nii0lil, ni1iOli}),
	.o(wire_nl111ii_o),
	.sel({(~ n0OiO), n0OiO, 1'b0}));
	defparam
		nl111ii.width_data = 3,
		nl111ii.width_sel = 3;
	oper_selector   nl111il
	( 
	.data({1'b0, nii0lli, ni1iOli}),
	.o(wire_nl111il_o),
	.sel({(~ n0OiO), n0OiO, 1'b0}));
	defparam
		nl111il.width_data = 3,
		nl111il.width_sel = 3;
	oper_selector   nl111Ol
	( 
	.data({1'b1, (~ nli11lO), nl00lli, {15{1'b0}}}),
	.o(wire_nl111Ol_o),
	.sel({ni1010l, ni1010i, ni1011O, {13{1'b0}}, ni1011l, (~ (((ni1010l | ni1010i) | ni1011O) | ni1011l))}));
	defparam
		nl111Ol.width_data = 18,
		nl111Ol.width_sel = 18;
	oper_selector   nl11Oii
	( 
	.data({1'b0, nil1i1O, ni1iOli}),
	.o(wire_nl11Oii_o),
	.sel({(~ n0Oil), n0Oil, 1'b0}));
	defparam
		nl11Oii.width_data = 3,
		nl11Oii.width_sel = 3;
	oper_selector   nl11Oil
	( 
	.data({1'b0, nil1i0i, ni1iOli}),
	.o(wire_nl11Oil_o),
	.sel({(~ n0Oil), n0Oil, 1'b0}));
	defparam
		nl11Oil.width_data = 3,
		nl11Oil.width_sel = 3;
	oper_selector   nl11OiO
	( 
	.data({1'b0, nil1i0l, ni1iOli}),
	.o(wire_nl11OiO_o),
	.sel({(~ n0Oil), n0Oil, 1'b0}));
	defparam
		nl11OiO.width_data = 3,
		nl11OiO.width_sel = 3;
	oper_selector   nl11Oli
	( 
	.data({1'b0, nil1i0O, ni1iOli}),
	.o(wire_nl11Oli_o),
	.sel({(~ n0Oil), n0Oil, 1'b0}));
	defparam
		nl11Oli.width_data = 3,
		nl11Oli.width_sel = 3;
	oper_selector   nl11Oll
	( 
	.data({1'b0, nil1iii, ni1iOli}),
	.o(wire_nl11Oll_o),
	.sel({(~ n0Oil), n0Oil, 1'b0}));
	defparam
		nl11Oll.width_data = 3,
		nl11Oll.width_sel = 3;
	oper_selector   nl11OlO
	( 
	.data({1'b0, nil1iil, ni1iOli}),
	.o(wire_nl11OlO_o),
	.sel({(~ n0Oil), n0Oil, 1'b0}));
	defparam
		nl11OlO.width_data = 3,
		nl11OlO.width_sel = 3;
	oper_selector   nl11OOi
	( 
	.data({1'b0, nil1iiO, ni1iOli}),
	.o(wire_nl11OOi_o),
	.sel({(~ n0Oil), n0Oil, 1'b0}));
	defparam
		nl11OOi.width_data = 3,
		nl11OOi.width_sel = 3;
	oper_selector   nl11OOl
	( 
	.data({1'b0, nil1ili, ni1iOli}),
	.o(wire_nl11OOl_o),
	.sel({(~ n0Oil), n0Oil, 1'b0}));
	defparam
		nl11OOl.width_data = 3,
		nl11OOl.width_sel = 3;
	oper_selector   nl11OOO
	( 
	.data({1'b0, nil1ill, ni1iOli}),
	.o(wire_nl11OOO_o),
	.sel({(~ n0Oil), n0Oil, 1'b0}));
	defparam
		nl11OOO.width_data = 3,
		nl11OOO.width_sel = 3;
	oper_selector   nl1l0lO
	( 
	.data({1'b1, nilOl0l, ni1iOli}),
	.o(wire_nl1l0lO_o),
	.sel({(~ n00il), n00il, 1'b0}));
	defparam
		nl1l0lO.width_data = 3,
		nl1l0lO.width_sel = 3;
	oper_selector   nl1l0Oi
	( 
	.data({1'b1, nilOl0O, ni1iOli}),
	.o(wire_nl1l0Oi_o),
	.sel({(~ n00il), n00il, 1'b0}));
	defparam
		nl1l0Oi.width_data = 3,
		nl1l0Oi.width_sel = 3;
	oper_selector   nl1l0Ol
	( 
	.data({1'b1, nilOlii, ni1iOli}),
	.o(wire_nl1l0Ol_o),
	.sel({(~ n00il), n00il, 1'b0}));
	defparam
		nl1l0Ol.width_data = 3,
		nl1l0Ol.width_sel = 3;
	oper_selector   nl1l0OO
	( 
	.data({1'b1, nilOlil, ni1iOli}),
	.o(wire_nl1l0OO_o),
	.sel({(~ n00il), n00il, 1'b0}));
	defparam
		nl1l0OO.width_data = 3,
		nl1l0OO.width_sel = 3;
	oper_selector   nl1li0i
	( 
	.data({1'b1, nilOlOi, ni1iOli}),
	.o(wire_nl1li0i_o),
	.sel({(~ n00il), n00il, 1'b0}));
	defparam
		nl1li0i.width_data = 3,
		nl1li0i.width_sel = 3;
	oper_selector   nl1li1i
	( 
	.data({1'b1, nilOliO, ni1iOli}),
	.o(wire_nl1li1i_o),
	.sel({(~ n00il), n00il, 1'b0}));
	defparam
		nl1li1i.width_data = 3,
		nl1li1i.width_sel = 3;
	oper_selector   nl1li1l
	( 
	.data({1'b1, nilOlli, ni1iOli}),
	.o(wire_nl1li1l_o),
	.sel({(~ n00il), n00il, 1'b0}));
	defparam
		nl1li1l.width_data = 3,
		nl1li1l.width_sel = 3;
	oper_selector   nl1li1O
	( 
	.data({1'b1, nilOlll, ni1iOli}),
	.o(wire_nl1li1O_o),
	.sel({(~ n00il), n00il, 1'b0}));
	defparam
		nl1li1O.width_data = 3,
		nl1li1O.width_sel = 3;
	oper_selector   nl1liOi
	( 
	.data({1'b0, nilOl0l, ni1iOli}),
	.o(wire_nl1liOi_o),
	.sel({(~ n0Oll), n0Oll, 1'b0}));
	defparam
		nl1liOi.width_data = 3,
		nl1liOi.width_sel = 3;
	oper_selector   nl1liOl
	( 
	.data({1'b0, nilOl0O, ni1iOli}),
	.o(wire_nl1liOl_o),
	.sel({(~ n0Oll), n0Oll, 1'b0}));
	defparam
		nl1liOl.width_data = 3,
		nl1liOl.width_sel = 3;
	oper_selector   nl1liOO
	( 
	.data({1'b0, nilOlii, ni1iOli}),
	.o(wire_nl1liOO_o),
	.sel({(~ n0Oll), n0Oll, 1'b0}));
	defparam
		nl1liOO.width_data = 3,
		nl1liOO.width_sel = 3;
	oper_selector   nl1ll0i
	( 
	.data({1'b0, nilOlll, ni1iOli}),
	.o(wire_nl1ll0i_o),
	.sel({(~ n0Oll), n0Oll, 1'b0}));
	defparam
		nl1ll0i.width_data = 3,
		nl1ll0i.width_sel = 3;
	oper_selector   nl1ll0l
	( 
	.data({1'b0, nilOlOi, ni1iOli}),
	.o(wire_nl1ll0l_o),
	.sel({(~ n0Oll), n0Oll, 1'b0}));
	defparam
		nl1ll0l.width_data = 3,
		nl1ll0l.width_sel = 3;
	oper_selector   nl1ll1i
	( 
	.data({1'b0, nilOlil, ni1iOli}),
	.o(wire_nl1ll1i_o),
	.sel({(~ n0Oll), n0Oll, 1'b0}));
	defparam
		nl1ll1i.width_data = 3,
		nl1ll1i.width_sel = 3;
	oper_selector   nl1ll1l
	( 
	.data({1'b0, nilOliO, ni1iOli}),
	.o(wire_nl1ll1l_o),
	.sel({(~ n0Oll), n0Oll, 1'b0}));
	defparam
		nl1ll1l.width_data = 3,
		nl1ll1l.width_sel = 3;
	oper_selector   nl1ll1O
	( 
	.data({1'b0, nilOlli, ni1iOli}),
	.o(wire_nl1ll1O_o),
	.sel({(~ n0Oll), n0Oll, 1'b0}));
	defparam
		nl1ll1O.width_data = 3,
		nl1ll1O.width_sel = 3;
	oper_selector   nl1llii
	( 
	.data({1'b1, (ni1iiOl | ((~ (nl1i0Oi & nli100O)) & nli101O)), ni1iOli}),
	.o(wire_nl1llii_o),
	.sel({(~ n0Oll), n0Oll, 1'b0}));
	defparam
		nl1llii.width_data = 3,
		nl1llii.width_sel = 3;
	oper_selector   nl1lliO
	( 
	.data({ni1iiOl, (~ (nl1i0OO | nl1i0Oi)), ni1iOli}),
	.o(wire_nl1lliO_o),
	.sel({(~ n00il), n00il, 1'b0}));
	defparam
		nl1lliO.width_data = 3,
		nl1lliO.width_sel = 3;
	assign
		alpha_in_0_ready = nilOi0l,
		alpha_in_1_ready = niO00lO,
		control_av_readdata = {wire_niOl0il_q_b[15:0]},
		din_0_ready = nil101O,
		din_1_ready = nilO00l,
		dout_data = {niOiO0l, niOiO1O, niOiO1l, niOiO1i, niOilOO, niOilOl, niOilOi, niOillO, niOilll, niOilli, niOiliO, niOilil, niOilii, niOil0O, niOil0l, niOil0i, niOil1O, niOil1l, niOil1i, niOiiOO, niOiiOl, niOiiOi, niOiilO, niOiill},
		dout_endofpacket = niOii1l,
		dout_startofpacket = niOii0i,
		dout_valid = niOiOii,
		n0OOili = ((((~ n00ii) & (~ n000O)) & n000l) & (~ n000i)),
		n0OOill = ((((~ n00ii) & (~ n000O)) & n000l) & n000i),
		n0OOilO = ((((~ n00ii) & n000O) & (~ n000l)) & (~ n000i)),
		n0OOiOi = ((((~ n00ii) & n000O) & (~ n000l)) & n000i),
		n0OOiOl = (((n00ii & (~ n000O)) & (~ n000l)) & (~ n000i)),
		n0OOiOO = (((n00ii & (~ n000O)) & (~ n000l)) & n000i),
		n0OOl0i = (((~ n0lil) & (~ n0lii)) & n0l0O),
		n0OOl0l = (((~ n10ll) & (~ n10li)) & (~ n10iO)),
		n0OOl0O = ((n10ll & (~ n10li)) & (~ n10iO)),
		n0OOl1i = (((~ n0lil) & (~ n0lii)) & (~ n0l0O)),
		n0OOl1l = ((n0lil & (~ n0lii)) & (~ n0l0O)),
		n0OOl1O = (((~ n0lil) & n0lii) & (~ n0l0O)),
		n0OOlii = (((~ n10ll) & n10li) & (~ n10iO)),
		n0OOlil = (((~ n10ll) & (~ n10li)) & n10iO),
		n0OOliO = (n0OOO0O & ((~ n0OOOii) | n0OOOil)),
		n0OOlli = ((~ n0OOO0O) & (n0OOOii & (~ n0OOOil))),
		n0OOlll = (n0OOO0O & (n0OOOil | (~ ni0101l))),
		n0OOllO = ((~ n0OOO0O) & ((~ n0OOOil) & ni0101l)),
		n0OOlOi = (n0OOO0O & (n0OOOil | (~ ni01lil))),
		n0OOlOl = ((~ n0OOO0O) & ((~ n0OOOil) & ni01lil)),
		n0OOlOO = (n0OOO0O & ((n0OOO0l & (ni01lli & ni01liO)) | ((~ n0OOO0l) & n0OOO1l))),
		n0OOO0i = ((~ ni01lli) & ni01liO),
		n0OOO0l = ((~ n0OOOil) & ni01lil),
		n0OOO0O = (((~ ni1iili) & wire_ni011ii_o) & (~ ni01iil)),
		n0OOO1i = (n0OOO0O & ((n0OOO0l & n0OOO1l) | ((~ n0OOO0l) & n0OOO0i))),
		n0OOO1l = (ni01lli & (~ ni01liO)),
		n0OOO1O = (n0OOO0O & ((n0OOO0l & n0OOO0i) | ((~ n0OOO0l) & ((~ ni01lli) & (~ ni01liO))))),
		n0OOOii = (((wire_nii111l_o | n0OOOiO) & (~ ni0100O)) & (~ n0OOOil)),
		n0OOOil = ((~ ((~ ni1iiii) & ni0Oi0l)) & ni0Oi0i),
		n0OOOiO = ((~ ni1iiii) & wire_ni011Ol_o),
		n0OOOli = (((~ n11ll) & (~ n11iO)) & (~ n11il)),
		n0OOOll = ((n11ll & (~ n11iO)) & (~ n11il)),
		n0OOOlO = (((~ n11ll) & n11iO) & (~ n11il)),
		n0OOOOi = (((~ n11ll) & (~ n11iO)) & n11il),
		n0OOOOl = ((~ ni1iiii) & wire_nii11iO_o),
		n0OOOOO = (n10Oi & ((~ ni1iiii) & nl0li0i)),
		ni1000i = (n00ll & (~ ni1iili)),
		ni1000l = (n1ill & (~ ni1iili)),
		ni1000O = (n1ill & (~ ni1iili)),
		ni1001i = (n01Oi & (~ ni1iili)),
		ni1001l = (n00ll & (~ ni1iili)),
		ni1001O = (n00ll & (~ ni1iili)),
		ni100ii = (n1ill & (~ ni1iili)),
		ni100il = (n01iO & ((~ ni1iili) & wire_nl1llii_o)),
		ni100iO = (n010O & (~ ni1iili)),
		ni100li = (n010O & (~ ni1iili)),
		ni100ll = (nlOOOi & (~ ni1iiii)),
		ni100lO = (nlO10l & (~ ni1iiii)),
		ni100Oi = (nlOOOl & (~ ni1iiii)),
		ni100Ol = ((((((((((((((ni10iOl | ni10iOi) | ni10ilO) | ni10ill) | ni10ili) | ni10iiO) | ni10iil) | ni10iii) | ni10i0O) | ni10i0l) | ni10i0i) | ni10i1O) | ni10i1l) | ni10i1i) | ni100OO),
		ni100OO = ((((((((((((((~ n0l0l) & (~ n0l0i)) & (~ n0l1O)) & (~ n0l1l)) & (~ n0l1i)) & (~ n0iOO)) & (~ n0iOl)) & (~ n0iOi)) & (~ n0ilO)) & (~ n0ill)) & (~ n0ili)) & (~ n0iiO)) & (~ n0iil)) & (~ n0iii)),
		ni1010i = ((n0lii & (~ n00ii)) & (~ n000O)),
		ni1010l = (((~ n0lii) & (~ n00ii)) & n000O),
		ni1010O = (n0O1l & ((~ ni1iili) & wire_nl111Ol_o)),
		ni1011i = ((~ ni1iili) & wire_niOO0iO_o),
		ni1011l = (((~ n0lii) & (~ n00ii)) & (~ n000O)),
		ni1011O = (((~ n0lii) & n00ii) & (~ n000O)),
		ni101ii = (((~ n0lil) & (~ n01lO)) & (~ n01ll)),
		ni101il = (((~ n0lil) & n01lO) & (~ n01ll)),
		ni101iO = ((n0lil & (~ n01lO)) & (~ n01ll)),
		ni101li = (((~ n0lil) & (~ n01lO)) & n01ll),
		ni101ll = (n0lOl & ((~ ni1iili) & wire_nl1000O_o)),
		ni101lO = (n0O1i & ((~ ni1iili) & nl0l0Oi)),
		ni101Oi = (n0lOi & ((~ ni1iili) & nl0l0Oi)),
		ni101Ol = (n0lOO & ((~ ni1iili) & nl0l0Oi)),
		ni101OO = (n0llO & ((~ ni1iili) & nl0l0Oi)),
		ni10i0i = ((((((((((((((~ n0l0l) & (~ n0l0i)) & (~ n0l1O)) & n0l1l) & (~ n0l1i)) & (~ n0iOO)) & (~ n0iOl)) & (~ n0iOi)) & (~ n0ilO)) & (~ n0ill)) & (~ n0ili)) & (~ n0iiO)) & (~ n0iil)) & (~ n0iii)),
		ni10i0l = ((((((((((((((~ n0l0l) & (~ n0l0i)) & (~ n0l1O)) & (~ n0l1l)) & n0l1i) & (~ n0iOO)) & (~ n0iOl)) & (~ n0iOi)) & (~ n0ilO)) & (~ n0ill)) & (~ n0ili)) & (~ n0iiO)) & (~ n0iil)) & (~ n0iii)),
		ni10i0O = ((((((((((((((~ n0l0l) & (~ n0l0i)) & (~ n0l1O)) & (~ n0l1l)) & (~ n0l1i)) & n0iOO) & (~ n0iOl)) & (~ n0iOi)) & (~ n0ilO)) & (~ n0ill)) & (~ n0ili)) & (~ n0iiO)) & (~ n0iil)) & (~ n0iii)),
		ni10i1i = (((((((((((((n0l0l & (~ n0l0i)) & (~ n0l1O)) & (~ n0l1l)) & (~ n0l1i)) & (~ n0iOO)) & (~ n0iOl)) & (~ n0iOi)) & (~ n0ilO)) & (~ n0ill)) & (~ n0ili)) & (~ n0iiO)) & (~ n0iil)) & (~ n0iii)),
		ni10i1l = ((((((((((((((~ n0l0l) & n0l0i) & (~ n0l1O)) & (~ n0l1l)) & (~ n0l1i)) & (~ n0iOO)) & (~ n0iOl)) & (~ n0iOi)) & (~ n0ilO)) & (~ n0ill)) & (~ n0ili)) & (~ n0iiO)) & (~ n0iil)) & (~ n0iii)),
		ni10i1O = ((((((((((((((~ n0l0l) & (~ n0l0i)) & n0l1O) & (~ n0l1l)) & (~ n0l1i)) & (~ n0iOO)) & (~ n0iOl)) & (~ n0iOi)) & (~ n0ilO)) & (~ n0ill)) & (~ n0ili)) & (~ n0iiO)) & (~ n0iil)) & (~ n0iii)),
		ni10iii = ((((((((((((((~ n0l0l) & (~ n0l0i)) & (~ n0l1O)) & (~ n0l1l)) & (~ n0l1i)) & (~ n0iOO)) & n0iOl) & (~ n0iOi)) & (~ n0ilO)) & (~ n0ill)) & (~ n0ili)) & (~ n0iiO)) & (~ n0iil)) & (~ n0iii)),
		ni10iil = ((((((((((((((~ n0l0l) & (~ n0l0i)) & (~ n0l1O)) & (~ n0l1l)) & (~ n0l1i)) & (~ n0iOO)) & (~ n0iOl)) & n0iOi) & (~ n0ilO)) & (~ n0ill)) & (~ n0ili)) & (~ n0iiO)) & (~ n0iil)) & (~ n0iii)),
		ni10iiO = ((((((((((((((~ n0l0l) & (~ n0l0i)) & (~ n0l1O)) & (~ n0l1l)) & (~ n0l1i)) & (~ n0iOO)) & (~ n0iOl)) & (~ n0iOi)) & n0ilO) & (~ n0ill)) & (~ n0ili)) & (~ n0iiO)) & (~ n0iil)) & (~ n0iii)),
		ni10ili = ((((((((((((((~ n0l0l) & (~ n0l0i)) & (~ n0l1O)) & (~ n0l1l)) & (~ n0l1i)) & (~ n0iOO)) & (~ n0iOl)) & (~ n0iOi)) & (~ n0ilO)) & n0ill) & (~ n0ili)) & (~ n0iiO)) & (~ n0iil)) & (~ n0iii)),
		ni10ill = ((((((((((((((~ n0l0l) & (~ n0l0i)) & (~ n0l1O)) & (~ n0l1l)) & (~ n0l1i)) & (~ n0iOO)) & (~ n0iOl)) & (~ n0iOi)) & (~ n0ilO)) & (~ n0ill)) & n0ili) & (~ n0iiO)) & (~ n0iil)) & (~ n0iii)),
		ni10ilO = ((((((((((((((~ n0l0l) & (~ n0l0i)) & (~ n0l1O)) & (~ n0l1l)) & (~ n0l1i)) & (~ n0iOO)) & (~ n0iOl)) & (~ n0iOi)) & (~ n0ilO)) & (~ n0ill)) & (~ n0ili)) & n0iiO) & (~ n0iil)) & (~ n0iii)),
		ni10iOi = ((((((((((((((~ n0l0l) & (~ n0l0i)) & (~ n0l1O)) & (~ n0l1l)) & (~ n0l1i)) & (~ n0iOO)) & (~ n0iOl)) & (~ n0iOi)) & (~ n0ilO)) & (~ n0ill)) & (~ n0ili)) & (~ n0iiO)) & n0iil) & (~ n0iii)),
		ni10iOl = ((((((((((((((~ n0l0l) & (~ n0l0i)) & (~ n0l1O)) & (~ n0l1l)) & (~ n0l1i)) & (~ n0iOO)) & (~ n0iOl)) & (~ n0iOi)) & (~ n0ilO)) & (~ n0ill)) & (~ n0ili)) & (~ n0iiO)) & (~ n0iil)) & n0iii),
		ni10iOO = (((((ni10l0O | ni10l0l) | ni10l0i) | ni10l1O) | ni10l1l) | ni10l1i),
		ni10l0i = (((((~ n0i0i) & (~ n0i1O)) & n0i1l) & (~ n0i1i)) & (~ n00OO)),
		ni10l0l = (((((~ n0i0i) & (~ n0i1O)) & (~ n0i1l)) & n0i1i) & (~ n00OO)),
		ni10l0O = (((((~ n0i0i) & (~ n0i1O)) & (~ n0i1l)) & (~ n0i1i)) & n00OO),
		ni10l1i = (((((~ n0i0i) & (~ n0i1O)) & (~ n0i1l)) & (~ n0i1i)) & (~ n00OO)),
		ni10l1l = ((((n0i0i & (~ n0i1O)) & (~ n0i1l)) & (~ n0i1i)) & (~ n00OO)),
		ni10l1O = (((((~ n0i0i) & n0i1O) & (~ n0i1l)) & (~ n0i1i)) & (~ n00OO)),
		ni10lii = ((((((((ni10O1i | ni10lOO) | ni10lOl) | ni10lOi) | ni10llO) | ni10lll) | ni10lli) | ni10liO) | ni10lil),
		ni10lil = ((((((((~ n10il) & (~ n10ii)) & (~ n100O)) & (~ n100l)) & (~ n100i)) & (~ n101O)) & (~ n101l)) & (~ n101i)),
		ni10liO = (((((((n10il & (~ n10ii)) & (~ n100O)) & (~ n100l)) & (~ n100i)) & (~ n101O)) & (~ n101l)) & (~ n101i)),
		ni10lli = ((((((((~ n10il) & n10ii) & (~ n100O)) & (~ n100l)) & (~ n100i)) & (~ n101O)) & (~ n101l)) & (~ n101i)),
		ni10lll = ((((((((~ n10il) & (~ n10ii)) & n100O) & (~ n100l)) & (~ n100i)) & (~ n101O)) & (~ n101l)) & (~ n101i)),
		ni10llO = ((((((((~ n10il) & (~ n10ii)) & (~ n100O)) & n100l) & (~ n100i)) & (~ n101O)) & (~ n101l)) & (~ n101i)),
		ni10lOi = ((((((((~ n10il) & (~ n10ii)) & (~ n100O)) & (~ n100l)) & n100i) & (~ n101O)) & (~ n101l)) & (~ n101i)),
		ni10lOl = ((((((((~ n10il) & (~ n10ii)) & (~ n100O)) & (~ n100l)) & (~ n100i)) & n101O) & (~ n101l)) & (~ n101i)),
		ni10lOO = ((((((((~ n10il) & (~ n10ii)) & (~ n100O)) & (~ n100l)) & (~ n100i)) & (~ n101O)) & n101l) & (~ n101i)),
		ni10O0i = (n00ii & (~ ni1iili)),
		ni10O0l = (n01lO & (~ ni1iili)),
		ni10O0O = (n00il & (~ ni1iili)),
		ni10O1i = ((((((((~ n10il) & (~ n10ii)) & (~ n100O)) & (~ n100l)) & (~ n100i)) & (~ n101O)) & (~ n101l)) & n101i),
		ni10O1l = 1'b0,
		ni10O1O = (n0Oli & (~ ni1iili)),
		ni10Oii = (n01il & (~ ni1iili)),
		ni10Oil = (n01ii & (~ ni1iili)),
		ni10OiO = (n11li & (~ ni1iiii)),
		ni10Oli = (nlOOOO & (~ ni1iiii)),
		ni10Oll = ((((~ nl00O1i) & (~ nl00lOl)) & (~ nl00lOi)) & (~ nl00llO)),
		ni10OlO = ((((~ nl00Oli) & (~ nl00Oil)) & (~ nl00Oii)) & (~ nl00O0O)),
		ni10OOi = ((((((((~ nl1lO0i) & (~ nl1lO1l)) & (~ nl1lO1i)) & (~ nl1llOO)) & (~ nl1llOl)) & (~ nl1llOi)) & (~ nl1lllO)) & (~ nl1llll)),
		ni10OOl = ((((((((((~ (niOlOlO ^ nl0iili)) & (~ (niOlO1l ^ nl0i0OO))) & (~ (niOlO1O ^ nl0ii1i))) & (~ (niOlO0i ^ nl0ii1l))) & (~ (niOlO0l ^ nl0ii1O))) & (~ (niOlO0O ^ nl0ii0i))) & (~ (niOlOii ^ nl0ii0l))) & (~ (niOlOil ^ nl0ii0O))) & (~ (niOlOiO ^ nl0iiii))) & (~ (niOlOli ^ nl0iiil))),
		ni10OOO = ((((((((~ (nl0i1Ol ^ nl0Olii)) & (~ (nl0i10O ^ nl0OiOl))) & (~ (nl0i1ii ^ nl0OiOO))) & (~ (nl0i1il ^ nl0Ol1i))) & (~ (nl0i1iO ^ nl0Ol1l))) & (~ (nl0i1li ^ nl0Ol1O))) & (~ (nl0i1ll ^ nl0Ol0i))) & (~ (nl0i1lO ^ nl0Ol0l))),
		ni1100i = ((((~ n00Ol) & n00Oi) & (~ n00lO)) & (~ n00ll)),
		ni1100l = ((((~ n00Ol) & (~ n00Oi)) & n00lO) & (~ n00ll)),
		ni1100O = ((((~ n00Ol) & (~ n00Oi)) & (~ n00lO)) & n00ll),
		ni1101i = ((((ni1100O | ni1100l) | ni1100i) | ni1101O) | ni1101l),
		ni1101l = ((((~ n00Ol) & (~ n00Oi)) & (~ n00lO)) & (~ n00ll)),
		ni1101O = (((n00Ol & (~ n00Oi)) & (~ n00lO)) & (~ n00ll)),
		ni110ii = (wire_nilO00i_dataout | wire_nilO01O_dataout),
		ni110il = (din_1_valid & ((ni110OO & nil1O1i) | ((~ ni110OO) & ni110li))),
		ni110iO = (din_1_valid & ((ni110OO & ni110li) | ((~ ni110OO) & ni110lO))),
		ni110li = ((~ nil1O1i) & nil1lOO),
		ni110ll = (din_1_valid & ((ni110OO & ni110lO) | ((~ ni110OO) & (~ nil1lOi)))),
		ni110lO = ((~ nil1lOO) & nil1lOi),
		ni110Oi = (din_1_valid & (~ ni110OO)),
		ni110Ol = ((~ din_1_valid) & ni110OO),
		ni110OO = (((~ ni1iili) & ((nilO01l | nilO01i) & nil1lOi)) & (~ ((~ nil0O1l) & nil01ll))),
		ni1110i = ((~ n0i0O) & (~ n0i0l)),
		ni1110l = (n0i0O & (~ n0i0l)),
		ni1110O = ((~ n0i0O) & n0i0l),
		ni1111i = (n10lO & ((~ ni1iiii) & nl0li0i)),
		ni1111l = (n0O0i & (~ ni1iili)),
		ni1111O = (n0Oll & (~ ni1iili)),
		ni111ii = (wire_nil101l_dataout | wire_nil101i_dataout),
		ni111il = (din_0_valid & ((ni111OO & nii0lOl) | ((~ ni111OO) & ni111li))),
		ni111iO = (din_0_valid & ((ni111OO & ni111li) | ((~ ni111OO) & ni111lO))),
		ni111li = ((~ nii0lOl) & nii0lOi),
		ni111ll = (din_0_valid & ((ni111OO & ni111lO) | ((~ ni111OO) & (~ nii0lll)))),
		ni111lO = ((~ nii0lOi) & nii0lll),
		ni111Oi = (din_0_valid & (~ ni111OO)),
		ni111Ol = ((~ din_0_valid) & ni111OO),
		ni111OO = (((~ ni1iili) & ((nil11OO | nil11Ol) & nii0lll)) & (~ ((~ niiilOO) & niii1iO))),
		ni11i0i = (((n00lO & (~ n00ll)) & (~ n00li)) & (~ n00iO)),
		ni11i0l = ((((~ n00lO) & n00ll) & (~ n00li)) & (~ n00iO)),
		ni11i0O = ((((~ n00lO) & (~ n00ll)) & (~ n00li)) & n00iO),
		ni11i1i = ((((ni11i0O | ni11i0l) | ni11i0i) | ni11i1O) | ni11i1l),
		ni11i1l = ((((~ n00lO) & (~ n00ll)) & (~ n00li)) & (~ n00iO)),
		ni11i1O = ((((~ n00lO) & (~ n00ll)) & n00li) & (~ n00iO)),
		ni11iii = (wire_niO00ll_dataout | wire_niO00li_dataout),
		ni11iil = (alpha_in_1_valid & ((ni11iOO & nilOO1l) | ((~ ni11iOO) & ni11ili))),
		ni11iiO = (alpha_in_1_valid & ((ni11iOO & ni11ili) | ((~ ni11iOO) & ni11ilO))),
		ni11ili = ((~ nilOO1l) & nilOO1i),
		ni11ill = (alpha_in_1_valid & ((ni11iOO & ni11ilO) | ((~ ni11iOO) & (~ nilOlOl)))),
		ni11ilO = ((~ nilOO1i) & nilOlOl),
		ni11iOi = (alpha_in_1_valid & (~ ni11iOO)),
		ni11iOl = ((~ alpha_in_1_valid) & ni11iOO),
		ni11iOO = (((~ ni1iili) & ((niO00iO | niO00il) & nilOlOl)) & (~ ((~ niO11OO) & nilOOll))),
		ni11l0i = (((~ n11li) & (~ n111l)) & n111i),
		ni11l0l = ((((ni11lli | ni11liO) | ni11lil) | ni11lii) | ni11l0O),
		ni11l0O = ((((~ n100i) & (~ n11OO)) & (~ n11Ol)) & (~ n11Oi)),
		ni11l1i = (((~ n11li) & (~ n111l)) & (~ n111i)),
		ni11l1l = (((~ n11li) & n111l) & (~ n111i)),
		ni11l1O = ((n11li & (~ n111l)) & (~ n111i)),
		ni11lii = ((((~ n100i) & n11OO) & (~ n11Ol)) & (~ n11Oi)),
		ni11lil = ((((~ n100i) & (~ n11OO)) & n11Ol) & (~ n11Oi)),
		ni11liO = (((n100i & (~ n11OO)) & (~ n11Ol)) & (~ n11Oi)),
		ni11lli = ((((~ n100i) & (~ n11OO)) & (~ n11Ol)) & n11Oi),
		ni11lll = ((((ni11O1i | ni11lOO) | ni11lOl) | ni11lOi) | ni11llO),
		ni11llO = ((((~ n100i) & (~ n11OO)) & (~ n11Ol)) & (~ n11lO)),
		ni11lOi = ((((~ n100i) & n11OO) & (~ n11Ol)) & (~ n11lO)),
		ni11lOl = ((((~ n100i) & (~ n11OO)) & n11Ol) & (~ n11lO)),
		ni11lOO = (((n100i & (~ n11OO)) & (~ n11Ol)) & (~ n11lO)),
		ni11O0i = (((~ n100i) & n101l) & (~ n110O)),
		ni11O0l = ((n100i & (~ n101l)) & (~ n110O)),
		ni11O0O = (ni11Oii & ni1iiiO),
		ni11O1i = ((((~ n100i) & (~ n11OO)) & (~ n11Ol)) & n11lO),
		ni11O1l = (((~ n100i) & (~ n101l)) & (~ n110O)),
		ni11O1O = (((~ n100i) & (~ n101l)) & n110O),
		ni11Oii = ((~ ni1iiii) & (n10OO & ni1iiil)),
		ni11Oil = ((~ n0OiO) & (~ n0Oil)),
		ni11OiO = ((~ n0OiO) & n0Oil),
		ni11Oli = (n0OiO & (~ n0Oil)),
		ni11Oll = ((~ ni1iili) & (n0Oii | niOl0Ol)),
		ni11OlO = (n0lll & (~ ni1iili)),
		ni11OOi = (n0O1O & (~ ni1iili)),
		ni11OOl = ((~ ni1iili) & wire_niOlOOl_o),
		ni11OOO = (n0lli & (~ ni1iili)),
		ni1i00i = (n010O & (~ ni1iili)),
		ni1i01l = (n010O & (~ ni1iili)),
		ni1i0ii = (n010O & (~ ni1iili)),
		ni1i0li = (n010O & (~ ni1iili)),
		ni1i0lO = (n010O & (~ ni1iili)),
		ni1i0OO = (n010O & (~ ni1iili)),
		ni1i10i = (((((((nl1lO0i & nl1lO1l) & nl1lO1i) & nl1llOO) & nl1llOl) & nl1llOi) & nl1lllO) & nl1llll),
		ni1i10l = (((((((((((((((((((((((((~ nii1iii) & (~ nii1i0l)) & (~ nii1i0i)) & (~ nii1i1O)) & (~ nii1i1l)) & (~ nii1i1i)) & (~ nii10OO)) & (~ nii10Ol)) & (~ nii10Oi)) & (~ nii10lO)) & (~ nii10ll)) & (~ nii10li)) & (~ nii10iO)) & (~ nii10il)) & (~ nii10ii)) & (~ nii100O)) & (~ nii100l)) & (~ nii100i)) & (~ nii101O)) & (~ nii101l)) & (~ nii101i)) & nii11OO) & nii11Ol) & nii11Oi) & nii11lO),
		ni1i11i = (n0O0i & (~ ni1iili)),
		ni1i11l = ((((((((((~ (niOlili ^ nl0iili)) & (~ (niOl0OO ^ nl0i0OO))) & (~ (niOli1i ^ nl0ii1i))) & (~ (niOli1l ^ nl0ii1l))) & (~ (niOli1O ^ nl0ii1O))) & (~ (niOli0i ^ nl0ii0i))) & (~ (niOli0l ^ nl0ii0l))) & (~ (niOli0O ^ nl0ii0O))) & (~ (niOliii ^ nl0iiii))) & (~ (niOliil ^ nl0iiil))),
		ni1i11O = ((((((((((~ (niOO1ll ^ nl0iili)) & (~ (niOO11i ^ nl0i0OO))) & (~ (niOO11l ^ nl0ii1i))) & (~ (niOO11O ^ nl0ii1l))) & (~ (niOO10i ^ nl0ii1O))) & (~ (niOO10l ^ nl0ii0i))) & (~ (niOO10O ^ nl0ii0l))) & (~ (niOO1ii ^ nl0ii0O))) & (~ (niOO1il ^ nl0iiii))) & (~ (niOO1iO ^ nl0iiil))),
		ni1i1il = ((((~ nii1OlO) & (~ nii1Oli)) & (~ nii1OiO)) & (~ nii1Oil)),
		ni1i1iO = (n0Oll & (~ ni1iili)),
		ni1i1lO = (n0Oll & (~ ni1iili)),
		ni1i1OO = (n0Oll & (~ ni1iili)),
		ni1ii0i = (n10OO & (~ ni1iiii)),
		ni1ii0l = (n10OO & (~ ni1iiii)),
		ni1ii0O = (n110O & (~ ni1iiii)),
		ni1ii1l = (n110O & (~ ni1iiii)),
		ni1iiii = (nlO1Oi | ((ni0Oi0l & (~ ni0Oi0i)) | ((~ ni1iiiO) & (wire_niOi00O_o | (n10OO & ni1iiil))))),
		ni1iiil = (wire_niO0i1l_o & wire_niO0ili_o),
		ni1iiiO = (niOiOii | (~ niOii0l)),
		ni1iili = (((((wire_ni011ii_o & ni01iil) | (nil11OO & (~ nii0lll))) | (nilO01l & (~ nil1lOi))) | (niO00iO & (~ nilOlOl))) | nllOOO),
		ni1iilO = (((nl0l1ll & nl0li0i) | (~ nl0li0i)) & (~ nii1O0i)),
		ni1iiOi = ((nl0l1ll & nl0li0i) | (~ nl0li0i)),
		ni1iiOl = ((nli101O & nli100O) & nl1i0Oi),
		ni1iiOO = ((~ wire_nl01Oli_o) & ((~ ni1iiii) | nl001li)),
		ni1il1i = 1'b1,
		ni1il1l = ((~ wire_nl01O1i_o) & ((~ ni1iili) | nl01O0l)),
		ni1iOli = 1'b0;
endmodule //alpha_mixer
//synopsys translate_on
//VALID FILE
