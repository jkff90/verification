`include "wishbone_uvc/wishbone_common.svh"
`include "wishbone_uvc/wishbone_transaction.svh"
`include "wishbone_uvc/wishbone_config.svh"
`include "wishbone_uvc/wishbone_adapter.svh"
`include "wishbone_uvc/wishbone_sequencer.svh"
`include "wishbone_uvc/wishbone_driver.svh"
`include "wishbone_uvc/wishbone_monitor.svh"
`include "wishbone_uvc/wishbone_agent.svh"
`include "wishbone_uvc/wishbone_sequence.svh"
