
`include "env_uvc/avlst_video_env_config.svh"
`include "env_uvc/avlst_video_env.svh"
