//=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-
//  This file <amba_axi4_coverage.svh> is a part of <Verification> project
//  Copyright (C) 2018  An Pham (anphambk@gmail.com)
//
//  This program is free software: you can redistribute it and/or modify
//  it under the terms of the GNU General Public License as published by
//  the Free Software Foundation, either version 3 of the License, or
//  (at your option) any later version.
//
//  This program is distributed in the hope that it will be useful,
//  but WITHOUT ANY WARRANTY; without even the implied warranty of
//  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
//  GNU General Public License for more details.
//
//  You should have received a copy of the GNU General Public License
//  along with this program.  If not, see <http://www.gnu.org/licenses/>.
//=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-

`ifndef __AMBA_AXI4_COVERAGE_SVH__
`define __AMBA_AXI4_COVERAGE_SVH__

//------------------------------------------------------------------------------
// CLASS: amba_axi4_coverage
//
// Coverage collector for amba_axi4 protocol
//------------------------------------------------------------------------------
class amba_axi4_coverage extends uvm_component;
    //--- attributes ---
    
    protected amba_axi4_transaction m_trans; // proctected transaction to sample
    protected amba_axi4_config cfg;
    
    //--- TLM ports/exports ---
    
    // object: analysis_export
    // Coverage collector's analysis_export.
    // This port should be connected to monitor's analysis_port in order to sample the transactions.
    uvm_analysis_imp #(amba_axi4_transaction, amba_axi4_coverage) analysis_export;
    
    //--- coverage ---
    covergroup cg_trans;
        option.per_instance = 1;
    endgroup : cg_trans
    
    //--- factory registration ---
    `uvm_component_utils(amba_axi4_coverage)
    
    //--- methods ---
    extern function new(string name="amba_axi4_coverage", uvm_component parent=null);
    extern virtual function void build_phase(uvm_phase phase);
    extern virtual function void write(amba_axi4_transaction trans);
endclass : amba_axi4_coverage

//------------------------------------------------------------------------------
// +Constructor: new
//------------------------------------------------------------------------------
function amba_axi4_coverage::new(string name="amba_axi4_coverage", uvm_component parent=null);
    super.new(name, parent);
    cg_trans = new();
endfunction : new

//------------------------------------------------------------------------------
// +Function: build_phase
//------------------------------------------------------------------------------
function void amba_axi4_coverage::build_phase(uvm_phase phase);
    assert(uvm_config_db #(amba_axi4_config)::get(this, "", "cfg", cfg));
    analysis_export = new("analysis_export", this);
    super.build_phase(phase);
endfunction : build_phase

//------------------------------------------------------------------------------
// +Function: write
//------------------------------------------------------------------------------
function void amba_axi4_coverage::write(amba_axi4_transaction trans);
    m_trans = trans;
    cg_trans.sample();
endfunction : write

`endif /* __AMBA_AXI4_COVERAGE_SVH__ */
